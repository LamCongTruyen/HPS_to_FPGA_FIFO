// Copyright (C) 2025  Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Altera and sold by Altera or its authorized distributors.  Please
// refer to the Altera Software License Subscription Agreements 
// on the Quartus Prime software download page.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 24.1std.0 Build 1077 03/04/2025 SC Lite Edition"

// DATE "11/14/2025 00:07:06"

// 
// Device: Altera 5CSEMA5F31C6 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module Computer_System (
	clock_bridge_0_in_clk_clk,
	fifo_hps_to_fpga_out_readdata,
	fifo_hps_to_fpga_out_read,
	fifo_hps_to_fpga_out_waitrequest,
	fifo_hps_to_fpga_out_csr_address,
	fifo_hps_to_fpga_out_csr_read,
	fifo_hps_to_fpga_out_csr_writedata,
	fifo_hps_to_fpga_out_csr_write,
	fifo_hps_to_fpga_out_csr_readdata,
	hps_io_hps_io_emac1_inst_TX_CLK,
	hps_io_hps_io_emac1_inst_TXD0,
	hps_io_hps_io_emac1_inst_TXD1,
	hps_io_hps_io_emac1_inst_TXD2,
	hps_io_hps_io_emac1_inst_TXD3,
	hps_io_hps_io_emac1_inst_RXD0,
	hps_io_hps_io_emac1_inst_MDIO,
	hps_io_hps_io_emac1_inst_MDC,
	hps_io_hps_io_emac1_inst_RX_CTL,
	hps_io_hps_io_emac1_inst_TX_CTL,
	hps_io_hps_io_emac1_inst_RX_CLK,
	hps_io_hps_io_emac1_inst_RXD1,
	hps_io_hps_io_emac1_inst_RXD2,
	hps_io_hps_io_emac1_inst_RXD3,
	hps_io_hps_io_qspi_inst_IO0,
	hps_io_hps_io_qspi_inst_IO1,
	hps_io_hps_io_qspi_inst_IO2,
	hps_io_hps_io_qspi_inst_IO3,
	hps_io_hps_io_qspi_inst_SS0,
	hps_io_hps_io_qspi_inst_CLK,
	hps_io_hps_io_sdio_inst_CMD,
	hps_io_hps_io_sdio_inst_D0,
	hps_io_hps_io_sdio_inst_D1,
	hps_io_hps_io_sdio_inst_CLK,
	hps_io_hps_io_sdio_inst_D2,
	hps_io_hps_io_sdio_inst_D3,
	hps_io_hps_io_usb1_inst_D0,
	hps_io_hps_io_usb1_inst_D1,
	hps_io_hps_io_usb1_inst_D2,
	hps_io_hps_io_usb1_inst_D3,
	hps_io_hps_io_usb1_inst_D4,
	hps_io_hps_io_usb1_inst_D5,
	hps_io_hps_io_usb1_inst_D6,
	hps_io_hps_io_usb1_inst_D7,
	hps_io_hps_io_usb1_inst_CLK,
	hps_io_hps_io_usb1_inst_STP,
	hps_io_hps_io_usb1_inst_DIR,
	hps_io_hps_io_usb1_inst_NXT,
	hps_io_hps_io_spim1_inst_CLK,
	hps_io_hps_io_spim1_inst_MOSI,
	hps_io_hps_io_spim1_inst_MISO,
	hps_io_hps_io_spim1_inst_SS0,
	hps_io_hps_io_uart0_inst_RX,
	hps_io_hps_io_uart0_inst_TX,
	hps_io_hps_io_i2c0_inst_SDA,
	hps_io_hps_io_i2c0_inst_SCL,
	hps_io_hps_io_i2c1_inst_SDA,
	hps_io_hps_io_i2c1_inst_SCL,
	hps_io_hps_io_gpio_inst_GPIO09,
	hps_io_hps_io_gpio_inst_GPIO35,
	hps_io_hps_io_gpio_inst_GPIO40,
	hps_io_hps_io_gpio_inst_GPIO41,
	hps_io_hps_io_gpio_inst_GPIO48,
	hps_io_hps_io_gpio_inst_GPIO53,
	hps_io_hps_io_gpio_inst_GPIO54,
	hps_io_hps_io_gpio_inst_GPIO61,
	memory_mem_a,
	memory_mem_ba,
	memory_mem_ck,
	memory_mem_ck_n,
	memory_mem_cke,
	memory_mem_cs_n,
	memory_mem_ras_n,
	memory_mem_cas_n,
	memory_mem_we_n,
	memory_mem_reset_n,
	memory_mem_dq,
	memory_mem_dqs,
	memory_mem_dqs_n,
	memory_mem_odt,
	memory_mem_dm,
	memory_oct_rzqin,
	onchip_sram_s1_address,
	onchip_sram_s1_clken,
	onchip_sram_s1_chipselect,
	onchip_sram_s1_write,
	onchip_sram_s1_readdata,
	onchip_sram_s1_writedata,
	onchip_sram_s1_byteenable,
	sdram_clk_clk,
	system_pll_ref_clk_clk,
	system_pll_ref_reset_reset)/* synthesis synthesis_greybox=0 */;
input 	clock_bridge_0_in_clk_clk;
output 	[31:0] fifo_hps_to_fpga_out_readdata;
input 	fifo_hps_to_fpga_out_read;
output 	fifo_hps_to_fpga_out_waitrequest;
input 	[2:0] fifo_hps_to_fpga_out_csr_address;
input 	fifo_hps_to_fpga_out_csr_read;
input 	[31:0] fifo_hps_to_fpga_out_csr_writedata;
input 	fifo_hps_to_fpga_out_csr_write;
output 	[31:0] fifo_hps_to_fpga_out_csr_readdata;
output 	hps_io_hps_io_emac1_inst_TX_CLK;
output 	hps_io_hps_io_emac1_inst_TXD0;
output 	hps_io_hps_io_emac1_inst_TXD1;
output 	hps_io_hps_io_emac1_inst_TXD2;
output 	hps_io_hps_io_emac1_inst_TXD3;
input 	hps_io_hps_io_emac1_inst_RXD0;
inout 	hps_io_hps_io_emac1_inst_MDIO;
output 	hps_io_hps_io_emac1_inst_MDC;
input 	hps_io_hps_io_emac1_inst_RX_CTL;
output 	hps_io_hps_io_emac1_inst_TX_CTL;
input 	hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_io_hps_io_emac1_inst_RXD1;
input 	hps_io_hps_io_emac1_inst_RXD2;
input 	hps_io_hps_io_emac1_inst_RXD3;
inout 	hps_io_hps_io_qspi_inst_IO0;
inout 	hps_io_hps_io_qspi_inst_IO1;
inout 	hps_io_hps_io_qspi_inst_IO2;
inout 	hps_io_hps_io_qspi_inst_IO3;
output 	hps_io_hps_io_qspi_inst_SS0;
output 	hps_io_hps_io_qspi_inst_CLK;
inout 	hps_io_hps_io_sdio_inst_CMD;
inout 	hps_io_hps_io_sdio_inst_D0;
inout 	hps_io_hps_io_sdio_inst_D1;
output 	hps_io_hps_io_sdio_inst_CLK;
inout 	hps_io_hps_io_sdio_inst_D2;
inout 	hps_io_hps_io_sdio_inst_D3;
inout 	hps_io_hps_io_usb1_inst_D0;
inout 	hps_io_hps_io_usb1_inst_D1;
inout 	hps_io_hps_io_usb1_inst_D2;
inout 	hps_io_hps_io_usb1_inst_D3;
inout 	hps_io_hps_io_usb1_inst_D4;
inout 	hps_io_hps_io_usb1_inst_D5;
inout 	hps_io_hps_io_usb1_inst_D6;
inout 	hps_io_hps_io_usb1_inst_D7;
input 	hps_io_hps_io_usb1_inst_CLK;
output 	hps_io_hps_io_usb1_inst_STP;
input 	hps_io_hps_io_usb1_inst_DIR;
input 	hps_io_hps_io_usb1_inst_NXT;
output 	hps_io_hps_io_spim1_inst_CLK;
output 	hps_io_hps_io_spim1_inst_MOSI;
input 	hps_io_hps_io_spim1_inst_MISO;
output 	hps_io_hps_io_spim1_inst_SS0;
input 	hps_io_hps_io_uart0_inst_RX;
output 	hps_io_hps_io_uart0_inst_TX;
inout 	hps_io_hps_io_i2c0_inst_SDA;
inout 	hps_io_hps_io_i2c0_inst_SCL;
inout 	hps_io_hps_io_i2c1_inst_SDA;
inout 	hps_io_hps_io_i2c1_inst_SCL;
inout 	hps_io_hps_io_gpio_inst_GPIO09;
inout 	hps_io_hps_io_gpio_inst_GPIO35;
inout 	hps_io_hps_io_gpio_inst_GPIO40;
inout 	hps_io_hps_io_gpio_inst_GPIO41;
inout 	hps_io_hps_io_gpio_inst_GPIO48;
inout 	hps_io_hps_io_gpio_inst_GPIO53;
inout 	hps_io_hps_io_gpio_inst_GPIO54;
inout 	hps_io_hps_io_gpio_inst_GPIO61;
output 	[14:0] memory_mem_a;
output 	[2:0] memory_mem_ba;
output 	memory_mem_ck;
output 	memory_mem_ck_n;
output 	memory_mem_cke;
output 	memory_mem_cs_n;
output 	memory_mem_ras_n;
output 	memory_mem_cas_n;
output 	memory_mem_we_n;
output 	memory_mem_reset_n;
inout 	[31:0] memory_mem_dq;
inout 	[3:0] memory_mem_dqs;
inout 	[3:0] memory_mem_dqs_n;
output 	memory_mem_odt;
output 	[3:0] memory_mem_dm;
input 	memory_oct_rzqin;
input 	[7:0] onchip_sram_s1_address;
input 	onchip_sram_s1_clken;
input 	onchip_sram_s1_chipselect;
input 	onchip_sram_s1_write;
output 	[31:0] onchip_sram_s1_readdata;
input 	[31:0] onchip_sram_s1_writedata;
input 	[3:0] onchip_sram_s1_byteenable;
output 	sdram_clk_clk;
input 	system_pll_ref_clk_clk;
input 	system_pll_ref_reset_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arm_a9_hps|fpga_interfaces|h2f_rst_n[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARVALID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWVALID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_BREADY[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_RREADY[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WLAST[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WVALID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARBURST[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARBURST[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[6] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[7] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[8] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[9] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[10] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARID[11] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWBURST[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWBURST[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[6] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[7] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[8] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[9] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[10] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWID[11] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[6] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[7] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[8] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[9] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[10] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[11] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[12] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[13] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[14] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[15] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[16] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[17] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[18] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[19] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[20] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[21] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[22] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[23] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[24] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[25] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[26] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[27] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[28] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[29] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[30] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[31] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARVALID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWVALID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_BREADY[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_RREADY[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WLAST[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WVALID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARADDR[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARADDR[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARADDR[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARADDR[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARADDR[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARADDR[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARADDR[6] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARADDR[7] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARADDR[8] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARADDR[9] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARBURST[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARBURST[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARID[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARID[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARID[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARID[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARID[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARID[6] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARID[7] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARID[8] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARID[9] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARID[10] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARID[11] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARLEN[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARLEN[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARLEN[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARLEN[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARSIZE[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARSIZE[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_ARSIZE[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[6] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[7] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[8] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[9] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[10] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[11] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[12] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[13] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[14] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[15] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[16] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[17] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[18] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[19] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[20] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[21] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[22] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[23] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[24] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[25] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[26] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWADDR[27] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWBURST[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWBURST[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWID[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWID[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWID[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWID[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWID[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWID[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWID[6] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWID[7] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWID[8] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWID[9] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWID[10] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWID[11] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWLEN[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWLEN[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWLEN[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWLEN[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWSIZE[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWSIZE[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_AWSIZE[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[6] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[7] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[8] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[9] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[10] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[11] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[12] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[13] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[14] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[15] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[16] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[17] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[18] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[19] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[20] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[21] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[22] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[23] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[24] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[25] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[26] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[27] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[28] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[29] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[30] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[31] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[32] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[33] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[34] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[35] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[36] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[37] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[38] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[39] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[40] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[41] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[42] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[43] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[44] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[45] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[46] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[47] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[48] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[49] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[50] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[51] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[52] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[53] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[54] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[55] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[56] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[57] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[58] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[59] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[60] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[61] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[62] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[63] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[64] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[65] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[66] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[67] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[68] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[69] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[70] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[71] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[72] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[73] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[74] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[75] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[76] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[77] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[78] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[79] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[80] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[81] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[82] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[83] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[84] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[85] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[86] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[87] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[88] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[89] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[90] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[91] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[92] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[93] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[94] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[95] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[96] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[97] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[98] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[99] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[100] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[101] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[102] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[103] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[104] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[105] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[106] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[107] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[108] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[109] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[110] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[111] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[112] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[113] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[114] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[115] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[116] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[117] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[118] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[119] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[120] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[121] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[122] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[123] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[124] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[125] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[126] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WDATA[127] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[0] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[1] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[2] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[3] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[4] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[5] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[6] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[7] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[8] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[9] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[10] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[11] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[12] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[13] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[14] ;
wire \arm_a9_hps|fpga_interfaces|h2f_WSTRB[15] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[0] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[1] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[2] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[3] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[4] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[5] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[6] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[7] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[8] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[9] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[10] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[11] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[12] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[13] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[14] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[15] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[16] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[17] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[18] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[19] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[20] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[21] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[22] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[23] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[24] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[25] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[26] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[27] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[28] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[29] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[30] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[31] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[0] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[0] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[1] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[1] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[2] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[2] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[3] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[3] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[4] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[4] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[5] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[5] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[6] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[6] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[7] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[7] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[8] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[8] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[9] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[9] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[10] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[10] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[11] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[11] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[12] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[12] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[13] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[13] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[14] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[14] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[15] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[15] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[16] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[16] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[17] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[17] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[18] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[18] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[19] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[19] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[20] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[20] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[21] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[21] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[22] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[22] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[23] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[23] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[24] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[24] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[25] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[25] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[26] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[26] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[27] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[27] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[28] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[28] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[29] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[29] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[30] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[30] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_a[31] ;
wire \onchip_sram|the_altsyncram|auto_generated|q_b[31] ;
wire \system_pll|sys_pll|altera_pll_i|outclk_wire[1] ;
wire \system_pll|sys_pll|altera_pll_i|outclk_wire[0] ;
wire \system_pll|sys_pll|altera_pll_i|locked_wire[0] ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|op_2~13_sumout ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|op_2~25_sumout ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|op_2~29_sumout ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[5]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[6]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[7]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[8]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[9]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~combout ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[0]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[1]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[2]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[3]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[4]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[5]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[6]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[7]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_1|cmd_mux|sink1_ready~combout ;
wire \mm_interconnect_1|arm_a9_hps_h2f_lw_axi_master_agent|awready~0_combout ;
wire \mm_interconnect_1|rsp_demux|src0_valid~combout ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent|uncompressor|source_endofpacket~combout ;
wire \mm_interconnect_1|rsp_demux|src1_valid~0_combout ;
wire \mm_interconnect_1|arm_a9_hps_h2f_lw_axi_master_agent|wready~0_combout ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][88]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][89]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][90]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][91]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][92]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][93]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][94]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][95]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][96]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][97]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][98]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][99]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[0]~0_combout ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[1]~1_combout ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[2]~2_combout ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[3]~3_combout ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[4]~4_combout ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[5]~5_combout ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[6]~6_combout ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[7]~7_combout ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[34]~0_combout ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[32]~1_combout ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[33]~2_combout ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~4_combout ;
wire \mm_interconnect_0|cmd_mux_001|sink1_ready~combout ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~0_combout ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~1_combout ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~2_combout ;
wire \mm_interconnect_0|arm_a9_hps_h2f_axi_master_agent|awready~0_combout ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload[0]~combout ;
wire \mm_interconnect_0|rsp_mux_001|WideOr1~combout ;
wire \mm_interconnect_0|arm_a9_hps_h2f_axi_master_agent|wready~0_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[209]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[210]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[211]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[212]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[213]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[214]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[215]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[216]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[217]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[218]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[219]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[220]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[0]~1_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~4_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[2]~3_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[3]~5_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~6_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[5]~7_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~8_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[7]~9_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~10_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[9]~11_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[10]~13_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[11]~15_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[12]~17_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~12_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[14]~19_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[15]~21_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[16]~23_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~14_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[18]~25_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[19]~27_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~16_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[21]~29_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~18_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[23]~31_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~20_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[25]~33_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[26]~35_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[27]~37_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[28]~39_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~22_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[30]~41_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[31]~43_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[32]~45_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~26_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[34]~47_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[35]~49_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~28_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[37]~51_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~30_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[39]~53_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~32_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[41]~55_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[42]~57_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[43]~59_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[44]~61_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~34_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[46]~63_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[47]~65_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[48]~67_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~36_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[50]~69_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[51]~71_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~38_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[53]~73_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~40_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[55]~75_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~42_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[57]~77_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[58]~79_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[59]~81_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[60]~83_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~44_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[62]~85_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[63]~87_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[64]~89_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~48_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[66]~91_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[67]~93_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~50_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[69]~95_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~52_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[71]~97_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~54_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[73]~99_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[74]~101_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[75]~103_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[76]~105_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~56_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[78]~107_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[79]~109_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[80]~111_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~58_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[82]~113_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[83]~115_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~60_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[85]~117_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~62_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[87]~119_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~64_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[89]~121_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[90]~123_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[91]~125_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[92]~127_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~66_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[94]~129_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[95]~131_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[96]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~71_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[98]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[99]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~72_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[101]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~73_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[103]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~74_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[105]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[106]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[107]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[108]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~75_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[110]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[111]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[112]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~76_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[114]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[115]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~77_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[117]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~78_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[119]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~79_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[121]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[122]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[123]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[124]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~80_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[126]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[127]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[209]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[210]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[211]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[212]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[213]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[214]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[215]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[216]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[217]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[218]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[219]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[220]~combout ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_agent|m0_write~0_combout ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ;
wire \mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ;
wire \rst_controller|r_sync_rst~q ;
wire \mm_interconnect_0|onchip_sram_s2_agent|m0_write~0_combout ;
wire \rst_controller|r_early_rst~q ;
wire \rst_controller_001|r_early_rst~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ;
wire \mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ;
wire \rst_controller_001|r_sync_rst~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent|m0_write~combout ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent|m0_read~0_combout ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[0]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[1]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[2]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[3]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[4]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[5]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[6]~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[7]~q ;
wire \rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~4_combout ;
wire \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~5_combout ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ;
wire \mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ;
wire \rst_controller_001|merged_reset~0_combout ;
wire \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_CLK_TX ;
wire \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ;
wire \arm_a9_hps|hps_io|border|intermediate[0] ;
wire \arm_a9_hps|hps_io|border|intermediate[1] ;
wire \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ;
wire \arm_a9_hps|hps_io|border|emac1_inst~emac_phy_txd ;
wire \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ;
wire \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ;
wire \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ;
wire \arm_a9_hps|hps_io|border|qspi_inst~O_QSPI_SCLK ;
wire \arm_a9_hps|hps_io|border|intermediate[2] ;
wire \arm_a9_hps|hps_io|border|intermediate[4] ;
wire \arm_a9_hps|hps_io|border|intermediate[6] ;
wire \arm_a9_hps|hps_io|border|intermediate[8] ;
wire \arm_a9_hps|hps_io|border|intermediate[3] ;
wire \arm_a9_hps|hps_io|border|intermediate[5] ;
wire \arm_a9_hps|hps_io|border|intermediate[7] ;
wire \arm_a9_hps|hps_io|border|intermediate[9] ;
wire \arm_a9_hps|hps_io|border|qspi_inst~O_QSPI_SS_N0 ;
wire \arm_a9_hps|hps_io|border|sdio_inst~sdmmc_cclk ;
wire \arm_a9_hps|hps_io|border|intermediate[10] ;
wire \arm_a9_hps|hps_io|border|intermediate[11] ;
wire \arm_a9_hps|hps_io|border|intermediate[12] ;
wire \arm_a9_hps|hps_io|border|intermediate[14] ;
wire \arm_a9_hps|hps_io|border|intermediate[16] ;
wire \arm_a9_hps|hps_io|border|intermediate[18] ;
wire \arm_a9_hps|hps_io|border|intermediate[13] ;
wire \arm_a9_hps|hps_io|border|intermediate[15] ;
wire \arm_a9_hps|hps_io|border|intermediate[17] ;
wire \arm_a9_hps|hps_io|border|intermediate[19] ;
wire \arm_a9_hps|hps_io|border|usb1_inst~usb_ulpi_stp ;
wire \arm_a9_hps|hps_io|border|intermediate[20] ;
wire \arm_a9_hps|hps_io|border|intermediate[22] ;
wire \arm_a9_hps|hps_io|border|intermediate[24] ;
wire \arm_a9_hps|hps_io|border|intermediate[26] ;
wire \arm_a9_hps|hps_io|border|intermediate[28] ;
wire \arm_a9_hps|hps_io|border|intermediate[30] ;
wire \arm_a9_hps|hps_io|border|intermediate[32] ;
wire \arm_a9_hps|hps_io|border|intermediate[34] ;
wire \arm_a9_hps|hps_io|border|intermediate[21] ;
wire \arm_a9_hps|hps_io|border|intermediate[23] ;
wire \arm_a9_hps|hps_io|border|intermediate[25] ;
wire \arm_a9_hps|hps_io|border|intermediate[27] ;
wire \arm_a9_hps|hps_io|border|intermediate[29] ;
wire \arm_a9_hps|hps_io|border|intermediate[31] ;
wire \arm_a9_hps|hps_io|border|intermediate[33] ;
wire \arm_a9_hps|hps_io|border|intermediate[35] ;
wire \arm_a9_hps|hps_io|border|spim1_inst~O_SPI_MASTER_SCLK ;
wire \arm_a9_hps|hps_io|border|spim1_inst~O_SPI_MASTER_SS_0_N ;
wire \arm_a9_hps|hps_io|border|intermediate[36] ;
wire \arm_a9_hps|hps_io|border|intermediate[37] ;
wire \arm_a9_hps|hps_io|border|uart0_inst~uart_txd ;
wire \arm_a9_hps|hps_io|border|intermediate[39] ;
wire \arm_a9_hps|hps_io|border|intermediate[38] ;
wire \arm_a9_hps|hps_io|border|intermediate[41] ;
wire \arm_a9_hps|hps_io|border|intermediate[40] ;
wire \arm_a9_hps|hps_io|border|intermediate[42] ;
wire \arm_a9_hps|hps_io|border|intermediate[43] ;
wire \arm_a9_hps|hps_io|border|intermediate[44] ;
wire \arm_a9_hps|hps_io|border|intermediate[46] ;
wire \arm_a9_hps|hps_io|border|intermediate[48] ;
wire \arm_a9_hps|hps_io|border|intermediate[50] ;
wire \arm_a9_hps|hps_io|border|intermediate[52] ;
wire \arm_a9_hps|hps_io|border|intermediate[54] ;
wire \arm_a9_hps|hps_io|border|intermediate[45] ;
wire \arm_a9_hps|hps_io|border|intermediate[47] ;
wire \arm_a9_hps|hps_io|border|intermediate[49] ;
wire \arm_a9_hps|hps_io|border|intermediate[51] ;
wire \arm_a9_hps|hps_io|border|intermediate[53] ;
wire \arm_a9_hps|hps_io|border|intermediate[55] ;
wire \arm_a9_hps|hps_io|border|intermediate[56] ;
wire \arm_a9_hps|hps_io|border|intermediate[57] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~input_o ;
wire \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD0~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD1~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD2~input_o ;
wire \hps_io_hps_io_emac1_inst_RXD3~input_o ;
wire \hps_io_hps_io_emac1_inst_RX_CLK~input_o ;
wire \hps_io_hps_io_emac1_inst_RX_CTL~input_o ;
wire \hps_io_hps_io_spim1_inst_MISO~input_o ;
wire \hps_io_hps_io_uart0_inst_RX~input_o ;
wire \hps_io_hps_io_usb1_inst_CLK~input_o ;
wire \hps_io_hps_io_usb1_inst_DIR~input_o ;
wire \hps_io_hps_io_usb1_inst_NXT~input_o ;
wire \memory_oct_rzqin~input_o ;
wire \fifo_hps_to_fpga_out_read~input_o ;
wire \clock_bridge_0_in_clk_clk~input_o ;
wire \fifo_hps_to_fpga_out_csr_address[2]~input_o ;
wire \fifo_hps_to_fpga_out_csr_address[0]~input_o ;
wire \fifo_hps_to_fpga_out_csr_address[1]~input_o ;
wire \fifo_hps_to_fpga_out_csr_read~input_o ;
wire \onchip_sram_s1_chipselect~input_o ;
wire \onchip_sram_s1_write~input_o ;
wire \onchip_sram_s1_clken~input_o ;
wire \onchip_sram_s1_writedata[0]~input_o ;
wire \onchip_sram_s1_address[0]~input_o ;
wire \onchip_sram_s1_address[1]~input_o ;
wire \onchip_sram_s1_address[2]~input_o ;
wire \onchip_sram_s1_address[3]~input_o ;
wire \onchip_sram_s1_address[4]~input_o ;
wire \onchip_sram_s1_address[5]~input_o ;
wire \onchip_sram_s1_address[6]~input_o ;
wire \onchip_sram_s1_address[7]~input_o ;
wire \onchip_sram_s1_byteenable[0]~input_o ;
wire \onchip_sram_s1_writedata[1]~input_o ;
wire \onchip_sram_s1_writedata[2]~input_o ;
wire \onchip_sram_s1_writedata[3]~input_o ;
wire \onchip_sram_s1_writedata[4]~input_o ;
wire \onchip_sram_s1_writedata[5]~input_o ;
wire \onchip_sram_s1_writedata[6]~input_o ;
wire \onchip_sram_s1_writedata[7]~input_o ;
wire \onchip_sram_s1_writedata[8]~input_o ;
wire \onchip_sram_s1_byteenable[1]~input_o ;
wire \onchip_sram_s1_writedata[9]~input_o ;
wire \onchip_sram_s1_writedata[10]~input_o ;
wire \onchip_sram_s1_writedata[11]~input_o ;
wire \onchip_sram_s1_writedata[12]~input_o ;
wire \onchip_sram_s1_writedata[13]~input_o ;
wire \onchip_sram_s1_writedata[14]~input_o ;
wire \onchip_sram_s1_writedata[15]~input_o ;
wire \onchip_sram_s1_writedata[16]~input_o ;
wire \onchip_sram_s1_byteenable[2]~input_o ;
wire \onchip_sram_s1_writedata[17]~input_o ;
wire \onchip_sram_s1_writedata[18]~input_o ;
wire \onchip_sram_s1_writedata[19]~input_o ;
wire \onchip_sram_s1_writedata[20]~input_o ;
wire \onchip_sram_s1_writedata[21]~input_o ;
wire \onchip_sram_s1_writedata[22]~input_o ;
wire \onchip_sram_s1_writedata[23]~input_o ;
wire \onchip_sram_s1_writedata[24]~input_o ;
wire \onchip_sram_s1_byteenable[3]~input_o ;
wire \onchip_sram_s1_writedata[25]~input_o ;
wire \onchip_sram_s1_writedata[26]~input_o ;
wire \onchip_sram_s1_writedata[27]~input_o ;
wire \onchip_sram_s1_writedata[28]~input_o ;
wire \onchip_sram_s1_writedata[29]~input_o ;
wire \onchip_sram_s1_writedata[30]~input_o ;
wire \onchip_sram_s1_writedata[31]~input_o ;
wire \system_pll_ref_clk_clk~input_o ;
wire \system_pll_ref_reset_reset~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[0]~input_o ;
wire \fifo_hps_to_fpga_out_csr_write~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[7]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[1]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[13]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[19]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[26]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[27]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[28]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[29]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[30]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[31]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[20]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[21]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[22]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[23]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[24]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[25]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[8]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[9]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[10]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[11]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[12]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[14]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[15]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[16]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[17]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[18]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[2]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[3]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[4]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[5]~input_o ;
wire \fifo_hps_to_fpga_out_csr_writedata[6]~input_o ;


Computer_System_Computer_System_mm_interconnect_0 mm_interconnect_0(
	.h2f_ARVALID_0(\arm_a9_hps|fpga_interfaces|h2f_ARVALID[0] ),
	.h2f_AWVALID_0(\arm_a9_hps|fpga_interfaces|h2f_AWVALID[0] ),
	.h2f_BREADY_0(\arm_a9_hps|fpga_interfaces|h2f_BREADY[0] ),
	.h2f_RREADY_0(\arm_a9_hps|fpga_interfaces|h2f_RREADY[0] ),
	.h2f_WLAST_0(\arm_a9_hps|fpga_interfaces|h2f_WLAST[0] ),
	.h2f_WVALID_0(\arm_a9_hps|fpga_interfaces|h2f_WVALID[0] ),
	.h2f_ARADDR_0(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[0] ),
	.h2f_ARADDR_1(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[1] ),
	.h2f_ARADDR_2(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[2] ),
	.h2f_ARADDR_3(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[3] ),
	.h2f_ARADDR_4(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[4] ),
	.h2f_ARADDR_5(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[5] ),
	.h2f_ARADDR_6(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[6] ),
	.h2f_ARADDR_7(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[7] ),
	.h2f_ARADDR_8(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[8] ),
	.h2f_ARADDR_9(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[9] ),
	.h2f_ARBURST_0(\arm_a9_hps|fpga_interfaces|h2f_ARBURST[0] ),
	.h2f_ARBURST_1(\arm_a9_hps|fpga_interfaces|h2f_ARBURST[1] ),
	.h2f_ARID_0(\arm_a9_hps|fpga_interfaces|h2f_ARID[0] ),
	.h2f_ARID_1(\arm_a9_hps|fpga_interfaces|h2f_ARID[1] ),
	.h2f_ARID_2(\arm_a9_hps|fpga_interfaces|h2f_ARID[2] ),
	.h2f_ARID_3(\arm_a9_hps|fpga_interfaces|h2f_ARID[3] ),
	.h2f_ARID_4(\arm_a9_hps|fpga_interfaces|h2f_ARID[4] ),
	.h2f_ARID_5(\arm_a9_hps|fpga_interfaces|h2f_ARID[5] ),
	.h2f_ARID_6(\arm_a9_hps|fpga_interfaces|h2f_ARID[6] ),
	.h2f_ARID_7(\arm_a9_hps|fpga_interfaces|h2f_ARID[7] ),
	.h2f_ARID_8(\arm_a9_hps|fpga_interfaces|h2f_ARID[8] ),
	.h2f_ARID_9(\arm_a9_hps|fpga_interfaces|h2f_ARID[9] ),
	.h2f_ARID_10(\arm_a9_hps|fpga_interfaces|h2f_ARID[10] ),
	.h2f_ARID_11(\arm_a9_hps|fpga_interfaces|h2f_ARID[11] ),
	.h2f_ARLEN_0(\arm_a9_hps|fpga_interfaces|h2f_ARLEN[0] ),
	.h2f_ARLEN_1(\arm_a9_hps|fpga_interfaces|h2f_ARLEN[1] ),
	.h2f_ARLEN_2(\arm_a9_hps|fpga_interfaces|h2f_ARLEN[2] ),
	.h2f_ARLEN_3(\arm_a9_hps|fpga_interfaces|h2f_ARLEN[3] ),
	.h2f_ARSIZE_0(\arm_a9_hps|fpga_interfaces|h2f_ARSIZE[0] ),
	.h2f_ARSIZE_1(\arm_a9_hps|fpga_interfaces|h2f_ARSIZE[1] ),
	.h2f_ARSIZE_2(\arm_a9_hps|fpga_interfaces|h2f_ARSIZE[2] ),
	.h2f_AWADDR_0(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[0] ),
	.h2f_AWADDR_1(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[1] ),
	.h2f_AWADDR_2(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[2] ),
	.h2f_AWADDR_3(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[3] ),
	.h2f_AWADDR_4(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[4] ),
	.h2f_AWADDR_5(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[5] ),
	.h2f_AWADDR_6(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[6] ),
	.h2f_AWADDR_7(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[7] ),
	.h2f_AWADDR_8(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[8] ),
	.h2f_AWADDR_9(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[9] ),
	.h2f_AWADDR_10(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[10] ),
	.h2f_AWADDR_11(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[11] ),
	.h2f_AWADDR_12(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[12] ),
	.h2f_AWADDR_13(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[13] ),
	.h2f_AWADDR_14(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[14] ),
	.h2f_AWADDR_15(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[15] ),
	.h2f_AWADDR_16(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[16] ),
	.h2f_AWADDR_17(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[17] ),
	.h2f_AWADDR_18(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[18] ),
	.h2f_AWADDR_19(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[19] ),
	.h2f_AWADDR_20(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[20] ),
	.h2f_AWADDR_21(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[21] ),
	.h2f_AWADDR_22(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[22] ),
	.h2f_AWADDR_23(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[23] ),
	.h2f_AWADDR_24(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[24] ),
	.h2f_AWADDR_25(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[25] ),
	.h2f_AWADDR_26(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[26] ),
	.h2f_AWADDR_27(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[27] ),
	.h2f_AWBURST_0(\arm_a9_hps|fpga_interfaces|h2f_AWBURST[0] ),
	.h2f_AWBURST_1(\arm_a9_hps|fpga_interfaces|h2f_AWBURST[1] ),
	.h2f_AWID_0(\arm_a9_hps|fpga_interfaces|h2f_AWID[0] ),
	.h2f_AWID_1(\arm_a9_hps|fpga_interfaces|h2f_AWID[1] ),
	.h2f_AWID_2(\arm_a9_hps|fpga_interfaces|h2f_AWID[2] ),
	.h2f_AWID_3(\arm_a9_hps|fpga_interfaces|h2f_AWID[3] ),
	.h2f_AWID_4(\arm_a9_hps|fpga_interfaces|h2f_AWID[4] ),
	.h2f_AWID_5(\arm_a9_hps|fpga_interfaces|h2f_AWID[5] ),
	.h2f_AWID_6(\arm_a9_hps|fpga_interfaces|h2f_AWID[6] ),
	.h2f_AWID_7(\arm_a9_hps|fpga_interfaces|h2f_AWID[7] ),
	.h2f_AWID_8(\arm_a9_hps|fpga_interfaces|h2f_AWID[8] ),
	.h2f_AWID_9(\arm_a9_hps|fpga_interfaces|h2f_AWID[9] ),
	.h2f_AWID_10(\arm_a9_hps|fpga_interfaces|h2f_AWID[10] ),
	.h2f_AWID_11(\arm_a9_hps|fpga_interfaces|h2f_AWID[11] ),
	.h2f_AWLEN_0(\arm_a9_hps|fpga_interfaces|h2f_AWLEN[0] ),
	.h2f_AWLEN_1(\arm_a9_hps|fpga_interfaces|h2f_AWLEN[1] ),
	.h2f_AWLEN_2(\arm_a9_hps|fpga_interfaces|h2f_AWLEN[2] ),
	.h2f_AWLEN_3(\arm_a9_hps|fpga_interfaces|h2f_AWLEN[3] ),
	.h2f_AWSIZE_0(\arm_a9_hps|fpga_interfaces|h2f_AWSIZE[0] ),
	.h2f_AWSIZE_1(\arm_a9_hps|fpga_interfaces|h2f_AWSIZE[1] ),
	.h2f_AWSIZE_2(\arm_a9_hps|fpga_interfaces|h2f_AWSIZE[2] ),
	.h2f_WDATA_0(\arm_a9_hps|fpga_interfaces|h2f_WDATA[0] ),
	.h2f_WDATA_1(\arm_a9_hps|fpga_interfaces|h2f_WDATA[1] ),
	.h2f_WDATA_2(\arm_a9_hps|fpga_interfaces|h2f_WDATA[2] ),
	.h2f_WDATA_3(\arm_a9_hps|fpga_interfaces|h2f_WDATA[3] ),
	.h2f_WDATA_4(\arm_a9_hps|fpga_interfaces|h2f_WDATA[4] ),
	.h2f_WDATA_5(\arm_a9_hps|fpga_interfaces|h2f_WDATA[5] ),
	.h2f_WDATA_6(\arm_a9_hps|fpga_interfaces|h2f_WDATA[6] ),
	.h2f_WDATA_7(\arm_a9_hps|fpga_interfaces|h2f_WDATA[7] ),
	.h2f_WDATA_8(\arm_a9_hps|fpga_interfaces|h2f_WDATA[8] ),
	.h2f_WDATA_9(\arm_a9_hps|fpga_interfaces|h2f_WDATA[9] ),
	.h2f_WDATA_10(\arm_a9_hps|fpga_interfaces|h2f_WDATA[10] ),
	.h2f_WDATA_11(\arm_a9_hps|fpga_interfaces|h2f_WDATA[11] ),
	.h2f_WDATA_12(\arm_a9_hps|fpga_interfaces|h2f_WDATA[12] ),
	.h2f_WDATA_13(\arm_a9_hps|fpga_interfaces|h2f_WDATA[13] ),
	.h2f_WDATA_14(\arm_a9_hps|fpga_interfaces|h2f_WDATA[14] ),
	.h2f_WDATA_15(\arm_a9_hps|fpga_interfaces|h2f_WDATA[15] ),
	.h2f_WDATA_16(\arm_a9_hps|fpga_interfaces|h2f_WDATA[16] ),
	.h2f_WDATA_17(\arm_a9_hps|fpga_interfaces|h2f_WDATA[17] ),
	.h2f_WDATA_18(\arm_a9_hps|fpga_interfaces|h2f_WDATA[18] ),
	.h2f_WDATA_19(\arm_a9_hps|fpga_interfaces|h2f_WDATA[19] ),
	.h2f_WDATA_20(\arm_a9_hps|fpga_interfaces|h2f_WDATA[20] ),
	.h2f_WDATA_21(\arm_a9_hps|fpga_interfaces|h2f_WDATA[21] ),
	.h2f_WDATA_22(\arm_a9_hps|fpga_interfaces|h2f_WDATA[22] ),
	.h2f_WDATA_23(\arm_a9_hps|fpga_interfaces|h2f_WDATA[23] ),
	.h2f_WDATA_24(\arm_a9_hps|fpga_interfaces|h2f_WDATA[24] ),
	.h2f_WDATA_25(\arm_a9_hps|fpga_interfaces|h2f_WDATA[25] ),
	.h2f_WDATA_26(\arm_a9_hps|fpga_interfaces|h2f_WDATA[26] ),
	.h2f_WDATA_27(\arm_a9_hps|fpga_interfaces|h2f_WDATA[27] ),
	.h2f_WDATA_28(\arm_a9_hps|fpga_interfaces|h2f_WDATA[28] ),
	.h2f_WDATA_29(\arm_a9_hps|fpga_interfaces|h2f_WDATA[29] ),
	.h2f_WDATA_30(\arm_a9_hps|fpga_interfaces|h2f_WDATA[30] ),
	.h2f_WDATA_31(\arm_a9_hps|fpga_interfaces|h2f_WDATA[31] ),
	.h2f_WDATA_32(\arm_a9_hps|fpga_interfaces|h2f_WDATA[32] ),
	.h2f_WDATA_33(\arm_a9_hps|fpga_interfaces|h2f_WDATA[33] ),
	.h2f_WDATA_34(\arm_a9_hps|fpga_interfaces|h2f_WDATA[34] ),
	.h2f_WDATA_35(\arm_a9_hps|fpga_interfaces|h2f_WDATA[35] ),
	.h2f_WDATA_36(\arm_a9_hps|fpga_interfaces|h2f_WDATA[36] ),
	.h2f_WDATA_37(\arm_a9_hps|fpga_interfaces|h2f_WDATA[37] ),
	.h2f_WDATA_38(\arm_a9_hps|fpga_interfaces|h2f_WDATA[38] ),
	.h2f_WDATA_39(\arm_a9_hps|fpga_interfaces|h2f_WDATA[39] ),
	.h2f_WDATA_40(\arm_a9_hps|fpga_interfaces|h2f_WDATA[40] ),
	.h2f_WDATA_41(\arm_a9_hps|fpga_interfaces|h2f_WDATA[41] ),
	.h2f_WDATA_42(\arm_a9_hps|fpga_interfaces|h2f_WDATA[42] ),
	.h2f_WDATA_43(\arm_a9_hps|fpga_interfaces|h2f_WDATA[43] ),
	.h2f_WDATA_44(\arm_a9_hps|fpga_interfaces|h2f_WDATA[44] ),
	.h2f_WDATA_45(\arm_a9_hps|fpga_interfaces|h2f_WDATA[45] ),
	.h2f_WDATA_46(\arm_a9_hps|fpga_interfaces|h2f_WDATA[46] ),
	.h2f_WDATA_47(\arm_a9_hps|fpga_interfaces|h2f_WDATA[47] ),
	.h2f_WDATA_48(\arm_a9_hps|fpga_interfaces|h2f_WDATA[48] ),
	.h2f_WDATA_49(\arm_a9_hps|fpga_interfaces|h2f_WDATA[49] ),
	.h2f_WDATA_50(\arm_a9_hps|fpga_interfaces|h2f_WDATA[50] ),
	.h2f_WDATA_51(\arm_a9_hps|fpga_interfaces|h2f_WDATA[51] ),
	.h2f_WDATA_52(\arm_a9_hps|fpga_interfaces|h2f_WDATA[52] ),
	.h2f_WDATA_53(\arm_a9_hps|fpga_interfaces|h2f_WDATA[53] ),
	.h2f_WDATA_54(\arm_a9_hps|fpga_interfaces|h2f_WDATA[54] ),
	.h2f_WDATA_55(\arm_a9_hps|fpga_interfaces|h2f_WDATA[55] ),
	.h2f_WDATA_56(\arm_a9_hps|fpga_interfaces|h2f_WDATA[56] ),
	.h2f_WDATA_57(\arm_a9_hps|fpga_interfaces|h2f_WDATA[57] ),
	.h2f_WDATA_58(\arm_a9_hps|fpga_interfaces|h2f_WDATA[58] ),
	.h2f_WDATA_59(\arm_a9_hps|fpga_interfaces|h2f_WDATA[59] ),
	.h2f_WDATA_60(\arm_a9_hps|fpga_interfaces|h2f_WDATA[60] ),
	.h2f_WDATA_61(\arm_a9_hps|fpga_interfaces|h2f_WDATA[61] ),
	.h2f_WDATA_62(\arm_a9_hps|fpga_interfaces|h2f_WDATA[62] ),
	.h2f_WDATA_63(\arm_a9_hps|fpga_interfaces|h2f_WDATA[63] ),
	.h2f_WDATA_64(\arm_a9_hps|fpga_interfaces|h2f_WDATA[64] ),
	.h2f_WDATA_65(\arm_a9_hps|fpga_interfaces|h2f_WDATA[65] ),
	.h2f_WDATA_66(\arm_a9_hps|fpga_interfaces|h2f_WDATA[66] ),
	.h2f_WDATA_67(\arm_a9_hps|fpga_interfaces|h2f_WDATA[67] ),
	.h2f_WDATA_68(\arm_a9_hps|fpga_interfaces|h2f_WDATA[68] ),
	.h2f_WDATA_69(\arm_a9_hps|fpga_interfaces|h2f_WDATA[69] ),
	.h2f_WDATA_70(\arm_a9_hps|fpga_interfaces|h2f_WDATA[70] ),
	.h2f_WDATA_71(\arm_a9_hps|fpga_interfaces|h2f_WDATA[71] ),
	.h2f_WDATA_72(\arm_a9_hps|fpga_interfaces|h2f_WDATA[72] ),
	.h2f_WDATA_73(\arm_a9_hps|fpga_interfaces|h2f_WDATA[73] ),
	.h2f_WDATA_74(\arm_a9_hps|fpga_interfaces|h2f_WDATA[74] ),
	.h2f_WDATA_75(\arm_a9_hps|fpga_interfaces|h2f_WDATA[75] ),
	.h2f_WDATA_76(\arm_a9_hps|fpga_interfaces|h2f_WDATA[76] ),
	.h2f_WDATA_77(\arm_a9_hps|fpga_interfaces|h2f_WDATA[77] ),
	.h2f_WDATA_78(\arm_a9_hps|fpga_interfaces|h2f_WDATA[78] ),
	.h2f_WDATA_79(\arm_a9_hps|fpga_interfaces|h2f_WDATA[79] ),
	.h2f_WDATA_80(\arm_a9_hps|fpga_interfaces|h2f_WDATA[80] ),
	.h2f_WDATA_81(\arm_a9_hps|fpga_interfaces|h2f_WDATA[81] ),
	.h2f_WDATA_82(\arm_a9_hps|fpga_interfaces|h2f_WDATA[82] ),
	.h2f_WDATA_83(\arm_a9_hps|fpga_interfaces|h2f_WDATA[83] ),
	.h2f_WDATA_84(\arm_a9_hps|fpga_interfaces|h2f_WDATA[84] ),
	.h2f_WDATA_85(\arm_a9_hps|fpga_interfaces|h2f_WDATA[85] ),
	.h2f_WDATA_86(\arm_a9_hps|fpga_interfaces|h2f_WDATA[86] ),
	.h2f_WDATA_87(\arm_a9_hps|fpga_interfaces|h2f_WDATA[87] ),
	.h2f_WDATA_88(\arm_a9_hps|fpga_interfaces|h2f_WDATA[88] ),
	.h2f_WDATA_89(\arm_a9_hps|fpga_interfaces|h2f_WDATA[89] ),
	.h2f_WDATA_90(\arm_a9_hps|fpga_interfaces|h2f_WDATA[90] ),
	.h2f_WDATA_91(\arm_a9_hps|fpga_interfaces|h2f_WDATA[91] ),
	.h2f_WDATA_92(\arm_a9_hps|fpga_interfaces|h2f_WDATA[92] ),
	.h2f_WDATA_93(\arm_a9_hps|fpga_interfaces|h2f_WDATA[93] ),
	.h2f_WDATA_94(\arm_a9_hps|fpga_interfaces|h2f_WDATA[94] ),
	.h2f_WDATA_95(\arm_a9_hps|fpga_interfaces|h2f_WDATA[95] ),
	.h2f_WDATA_96(\arm_a9_hps|fpga_interfaces|h2f_WDATA[96] ),
	.h2f_WDATA_97(\arm_a9_hps|fpga_interfaces|h2f_WDATA[97] ),
	.h2f_WDATA_98(\arm_a9_hps|fpga_interfaces|h2f_WDATA[98] ),
	.h2f_WDATA_99(\arm_a9_hps|fpga_interfaces|h2f_WDATA[99] ),
	.h2f_WDATA_100(\arm_a9_hps|fpga_interfaces|h2f_WDATA[100] ),
	.h2f_WDATA_101(\arm_a9_hps|fpga_interfaces|h2f_WDATA[101] ),
	.h2f_WDATA_102(\arm_a9_hps|fpga_interfaces|h2f_WDATA[102] ),
	.h2f_WDATA_103(\arm_a9_hps|fpga_interfaces|h2f_WDATA[103] ),
	.h2f_WDATA_104(\arm_a9_hps|fpga_interfaces|h2f_WDATA[104] ),
	.h2f_WDATA_105(\arm_a9_hps|fpga_interfaces|h2f_WDATA[105] ),
	.h2f_WDATA_106(\arm_a9_hps|fpga_interfaces|h2f_WDATA[106] ),
	.h2f_WDATA_107(\arm_a9_hps|fpga_interfaces|h2f_WDATA[107] ),
	.h2f_WDATA_108(\arm_a9_hps|fpga_interfaces|h2f_WDATA[108] ),
	.h2f_WDATA_109(\arm_a9_hps|fpga_interfaces|h2f_WDATA[109] ),
	.h2f_WDATA_110(\arm_a9_hps|fpga_interfaces|h2f_WDATA[110] ),
	.h2f_WDATA_111(\arm_a9_hps|fpga_interfaces|h2f_WDATA[111] ),
	.h2f_WDATA_112(\arm_a9_hps|fpga_interfaces|h2f_WDATA[112] ),
	.h2f_WDATA_113(\arm_a9_hps|fpga_interfaces|h2f_WDATA[113] ),
	.h2f_WDATA_114(\arm_a9_hps|fpga_interfaces|h2f_WDATA[114] ),
	.h2f_WDATA_115(\arm_a9_hps|fpga_interfaces|h2f_WDATA[115] ),
	.h2f_WDATA_116(\arm_a9_hps|fpga_interfaces|h2f_WDATA[116] ),
	.h2f_WDATA_117(\arm_a9_hps|fpga_interfaces|h2f_WDATA[117] ),
	.h2f_WDATA_118(\arm_a9_hps|fpga_interfaces|h2f_WDATA[118] ),
	.h2f_WDATA_119(\arm_a9_hps|fpga_interfaces|h2f_WDATA[119] ),
	.h2f_WDATA_120(\arm_a9_hps|fpga_interfaces|h2f_WDATA[120] ),
	.h2f_WDATA_121(\arm_a9_hps|fpga_interfaces|h2f_WDATA[121] ),
	.h2f_WDATA_122(\arm_a9_hps|fpga_interfaces|h2f_WDATA[122] ),
	.h2f_WDATA_123(\arm_a9_hps|fpga_interfaces|h2f_WDATA[123] ),
	.h2f_WDATA_124(\arm_a9_hps|fpga_interfaces|h2f_WDATA[124] ),
	.h2f_WDATA_125(\arm_a9_hps|fpga_interfaces|h2f_WDATA[125] ),
	.h2f_WDATA_126(\arm_a9_hps|fpga_interfaces|h2f_WDATA[126] ),
	.h2f_WDATA_127(\arm_a9_hps|fpga_interfaces|h2f_WDATA[127] ),
	.h2f_WSTRB_0(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[0] ),
	.h2f_WSTRB_1(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[1] ),
	.h2f_WSTRB_2(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[2] ),
	.h2f_WSTRB_3(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[3] ),
	.h2f_WSTRB_4(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[4] ),
	.h2f_WSTRB_5(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[5] ),
	.h2f_WSTRB_6(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[6] ),
	.h2f_WSTRB_7(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[7] ),
	.h2f_WSTRB_8(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[8] ),
	.h2f_WSTRB_9(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[9] ),
	.h2f_WSTRB_10(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[10] ),
	.h2f_WSTRB_11(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[11] ),
	.h2f_WSTRB_12(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[12] ),
	.h2f_WSTRB_13(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[13] ),
	.h2f_WSTRB_14(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[14] ),
	.h2f_WSTRB_15(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[15] ),
	.q_b_0(\onchip_sram|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\onchip_sram|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_2(\onchip_sram|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\onchip_sram|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_4(\onchip_sram|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\onchip_sram|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_6(\onchip_sram|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_7(\onchip_sram|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_8(\onchip_sram|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_9(\onchip_sram|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_10(\onchip_sram|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_11(\onchip_sram|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_12(\onchip_sram|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_13(\onchip_sram|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_14(\onchip_sram|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_15(\onchip_sram|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_16(\onchip_sram|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_17(\onchip_sram|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_18(\onchip_sram|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_19(\onchip_sram|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_20(\onchip_sram|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_21(\onchip_sram|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_22(\onchip_sram|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_23(\onchip_sram|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_24(\onchip_sram|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_25(\onchip_sram|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_26(\onchip_sram|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_27(\onchip_sram|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_28(\onchip_sram|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_29(\onchip_sram|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_30(\onchip_sram|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_31(\onchip_sram|the_altsyncram|auto_generated|q_b[31] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.op_2(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|op_2~13_sumout ),
	.op_21(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|op_2~25_sumout ),
	.op_22(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|op_2~29_sumout ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_4(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ),
	.int_nxt_addr_reg_dly_5(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[5]~q ),
	.int_nxt_addr_reg_dly_6(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[6]~q ),
	.int_nxt_addr_reg_dly_7(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[7]~q ),
	.int_nxt_addr_reg_dly_8(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[8]~q ),
	.int_nxt_addr_reg_dly_9(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[9]~q ),
	.in_ready_hold(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.source0_data_34(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[34]~0_combout ),
	.source0_data_32(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[32]~1_combout ),
	.source0_data_33(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[33]~2_combout ),
	.source0_data_35(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~4_combout ),
	.sink1_ready(\mm_interconnect_0|cmd_mux_001|sink1_ready~combout ),
	.wrfull(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~0_combout ),
	.wrfull1(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~1_combout ),
	.wrfull2(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~2_combout ),
	.ARM_A9_HPS_h2f_axi_master_awready(\mm_interconnect_0|arm_a9_hps_h2f_axi_master_agent|awready~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.src_payload_0(\mm_interconnect_0|rsp_mux_001|src_payload[0]~combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.ARM_A9_HPS_h2f_axi_master_wready(\mm_interconnect_0|arm_a9_hps_h2f_axi_master_agent|wready~0_combout ),
	.src_data_209(\mm_interconnect_0|rsp_mux|src_data[209]~combout ),
	.src_data_210(\mm_interconnect_0|rsp_mux|src_data[210]~combout ),
	.src_data_211(\mm_interconnect_0|rsp_mux|src_data[211]~combout ),
	.src_data_212(\mm_interconnect_0|rsp_mux|src_data[212]~combout ),
	.src_data_213(\mm_interconnect_0|rsp_mux|src_data[213]~combout ),
	.src_data_214(\mm_interconnect_0|rsp_mux|src_data[214]~combout ),
	.src_data_215(\mm_interconnect_0|rsp_mux|src_data[215]~combout ),
	.src_data_216(\mm_interconnect_0|rsp_mux|src_data[216]~combout ),
	.src_data_217(\mm_interconnect_0|rsp_mux|src_data[217]~combout ),
	.src_data_218(\mm_interconnect_0|rsp_mux|src_data[218]~combout ),
	.src_data_219(\mm_interconnect_0|rsp_mux|src_data[219]~combout ),
	.src_data_220(\mm_interconnect_0|rsp_mux|src_data[220]~combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux_001|src_data[0]~1_combout ),
	.src_payload(\mm_interconnect_0|rsp_mux_001|src_payload~4_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux_001|src_data[2]~3_combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux_001|src_data[3]~5_combout ),
	.src_payload1(\mm_interconnect_0|rsp_mux_001|src_payload~6_combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux_001|src_data[5]~7_combout ),
	.src_payload2(\mm_interconnect_0|rsp_mux_001|src_payload~8_combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux_001|src_data[7]~9_combout ),
	.src_payload3(\mm_interconnect_0|rsp_mux_001|src_payload~10_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux_001|src_data[9]~11_combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux_001|src_data[10]~13_combout ),
	.src_data_11(\mm_interconnect_0|rsp_mux_001|src_data[11]~15_combout ),
	.src_data_12(\mm_interconnect_0|rsp_mux_001|src_data[12]~17_combout ),
	.src_payload4(\mm_interconnect_0|rsp_mux_001|src_payload~12_combout ),
	.src_data_14(\mm_interconnect_0|rsp_mux_001|src_data[14]~19_combout ),
	.src_data_15(\mm_interconnect_0|rsp_mux_001|src_data[15]~21_combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux_001|src_data[16]~23_combout ),
	.src_payload5(\mm_interconnect_0|rsp_mux_001|src_payload~14_combout ),
	.src_data_18(\mm_interconnect_0|rsp_mux_001|src_data[18]~25_combout ),
	.src_data_19(\mm_interconnect_0|rsp_mux_001|src_data[19]~27_combout ),
	.src_payload6(\mm_interconnect_0|rsp_mux_001|src_payload~16_combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux_001|src_data[21]~29_combout ),
	.src_payload7(\mm_interconnect_0|rsp_mux_001|src_payload~18_combout ),
	.src_data_23(\mm_interconnect_0|rsp_mux_001|src_data[23]~31_combout ),
	.src_payload8(\mm_interconnect_0|rsp_mux_001|src_payload~20_combout ),
	.src_data_25(\mm_interconnect_0|rsp_mux_001|src_data[25]~33_combout ),
	.src_data_26(\mm_interconnect_0|rsp_mux_001|src_data[26]~35_combout ),
	.src_data_27(\mm_interconnect_0|rsp_mux_001|src_data[27]~37_combout ),
	.src_data_28(\mm_interconnect_0|rsp_mux_001|src_data[28]~39_combout ),
	.src_payload9(\mm_interconnect_0|rsp_mux_001|src_payload~22_combout ),
	.src_data_30(\mm_interconnect_0|rsp_mux_001|src_data[30]~41_combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux_001|src_data[31]~43_combout ),
	.src_data_32(\mm_interconnect_0|rsp_mux_001|src_data[32]~45_combout ),
	.src_payload10(\mm_interconnect_0|rsp_mux_001|src_payload~26_combout ),
	.src_data_34(\mm_interconnect_0|rsp_mux_001|src_data[34]~47_combout ),
	.src_data_35(\mm_interconnect_0|rsp_mux_001|src_data[35]~49_combout ),
	.src_payload11(\mm_interconnect_0|rsp_mux_001|src_payload~28_combout ),
	.src_data_37(\mm_interconnect_0|rsp_mux_001|src_data[37]~51_combout ),
	.src_payload12(\mm_interconnect_0|rsp_mux_001|src_payload~30_combout ),
	.src_data_39(\mm_interconnect_0|rsp_mux_001|src_data[39]~53_combout ),
	.src_payload13(\mm_interconnect_0|rsp_mux_001|src_payload~32_combout ),
	.src_data_41(\mm_interconnect_0|rsp_mux_001|src_data[41]~55_combout ),
	.src_data_42(\mm_interconnect_0|rsp_mux_001|src_data[42]~57_combout ),
	.src_data_43(\mm_interconnect_0|rsp_mux_001|src_data[43]~59_combout ),
	.src_data_44(\mm_interconnect_0|rsp_mux_001|src_data[44]~61_combout ),
	.src_payload14(\mm_interconnect_0|rsp_mux_001|src_payload~34_combout ),
	.src_data_46(\mm_interconnect_0|rsp_mux_001|src_data[46]~63_combout ),
	.src_data_47(\mm_interconnect_0|rsp_mux_001|src_data[47]~65_combout ),
	.src_data_48(\mm_interconnect_0|rsp_mux_001|src_data[48]~67_combout ),
	.src_payload15(\mm_interconnect_0|rsp_mux_001|src_payload~36_combout ),
	.src_data_50(\mm_interconnect_0|rsp_mux_001|src_data[50]~69_combout ),
	.src_data_51(\mm_interconnect_0|rsp_mux_001|src_data[51]~71_combout ),
	.src_payload16(\mm_interconnect_0|rsp_mux_001|src_payload~38_combout ),
	.src_data_53(\mm_interconnect_0|rsp_mux_001|src_data[53]~73_combout ),
	.src_payload17(\mm_interconnect_0|rsp_mux_001|src_payload~40_combout ),
	.src_data_55(\mm_interconnect_0|rsp_mux_001|src_data[55]~75_combout ),
	.src_payload18(\mm_interconnect_0|rsp_mux_001|src_payload~42_combout ),
	.src_data_57(\mm_interconnect_0|rsp_mux_001|src_data[57]~77_combout ),
	.src_data_58(\mm_interconnect_0|rsp_mux_001|src_data[58]~79_combout ),
	.src_data_59(\mm_interconnect_0|rsp_mux_001|src_data[59]~81_combout ),
	.src_data_60(\mm_interconnect_0|rsp_mux_001|src_data[60]~83_combout ),
	.src_payload19(\mm_interconnect_0|rsp_mux_001|src_payload~44_combout ),
	.src_data_62(\mm_interconnect_0|rsp_mux_001|src_data[62]~85_combout ),
	.src_data_63(\mm_interconnect_0|rsp_mux_001|src_data[63]~87_combout ),
	.src_data_64(\mm_interconnect_0|rsp_mux_001|src_data[64]~89_combout ),
	.src_payload20(\mm_interconnect_0|rsp_mux_001|src_payload~48_combout ),
	.src_data_66(\mm_interconnect_0|rsp_mux_001|src_data[66]~91_combout ),
	.src_data_67(\mm_interconnect_0|rsp_mux_001|src_data[67]~93_combout ),
	.src_payload21(\mm_interconnect_0|rsp_mux_001|src_payload~50_combout ),
	.src_data_69(\mm_interconnect_0|rsp_mux_001|src_data[69]~95_combout ),
	.src_payload22(\mm_interconnect_0|rsp_mux_001|src_payload~52_combout ),
	.src_data_71(\mm_interconnect_0|rsp_mux_001|src_data[71]~97_combout ),
	.src_payload23(\mm_interconnect_0|rsp_mux_001|src_payload~54_combout ),
	.src_data_73(\mm_interconnect_0|rsp_mux_001|src_data[73]~99_combout ),
	.src_data_74(\mm_interconnect_0|rsp_mux_001|src_data[74]~101_combout ),
	.src_data_75(\mm_interconnect_0|rsp_mux_001|src_data[75]~103_combout ),
	.src_data_76(\mm_interconnect_0|rsp_mux_001|src_data[76]~105_combout ),
	.src_payload24(\mm_interconnect_0|rsp_mux_001|src_payload~56_combout ),
	.src_data_78(\mm_interconnect_0|rsp_mux_001|src_data[78]~107_combout ),
	.src_data_79(\mm_interconnect_0|rsp_mux_001|src_data[79]~109_combout ),
	.src_data_80(\mm_interconnect_0|rsp_mux_001|src_data[80]~111_combout ),
	.src_payload25(\mm_interconnect_0|rsp_mux_001|src_payload~58_combout ),
	.src_data_82(\mm_interconnect_0|rsp_mux_001|src_data[82]~113_combout ),
	.src_data_83(\mm_interconnect_0|rsp_mux_001|src_data[83]~115_combout ),
	.src_payload26(\mm_interconnect_0|rsp_mux_001|src_payload~60_combout ),
	.src_data_85(\mm_interconnect_0|rsp_mux_001|src_data[85]~117_combout ),
	.src_payload27(\mm_interconnect_0|rsp_mux_001|src_payload~62_combout ),
	.src_data_87(\mm_interconnect_0|rsp_mux_001|src_data[87]~119_combout ),
	.src_payload28(\mm_interconnect_0|rsp_mux_001|src_payload~64_combout ),
	.src_data_89(\mm_interconnect_0|rsp_mux_001|src_data[89]~121_combout ),
	.src_data_90(\mm_interconnect_0|rsp_mux_001|src_data[90]~123_combout ),
	.src_data_91(\mm_interconnect_0|rsp_mux_001|src_data[91]~125_combout ),
	.src_data_92(\mm_interconnect_0|rsp_mux_001|src_data[92]~127_combout ),
	.src_payload29(\mm_interconnect_0|rsp_mux_001|src_payload~66_combout ),
	.src_data_94(\mm_interconnect_0|rsp_mux_001|src_data[94]~129_combout ),
	.src_data_95(\mm_interconnect_0|rsp_mux_001|src_data[95]~131_combout ),
	.src_data_96(\mm_interconnect_0|rsp_mux_001|src_data[96]~combout ),
	.src_payload30(\mm_interconnect_0|rsp_mux_001|src_payload~71_combout ),
	.src_data_98(\mm_interconnect_0|rsp_mux_001|src_data[98]~combout ),
	.src_data_99(\mm_interconnect_0|rsp_mux_001|src_data[99]~combout ),
	.src_payload31(\mm_interconnect_0|rsp_mux_001|src_payload~72_combout ),
	.src_data_101(\mm_interconnect_0|rsp_mux_001|src_data[101]~combout ),
	.src_payload32(\mm_interconnect_0|rsp_mux_001|src_payload~73_combout ),
	.src_data_103(\mm_interconnect_0|rsp_mux_001|src_data[103]~combout ),
	.src_payload33(\mm_interconnect_0|rsp_mux_001|src_payload~74_combout ),
	.src_data_105(\mm_interconnect_0|rsp_mux_001|src_data[105]~combout ),
	.src_data_106(\mm_interconnect_0|rsp_mux_001|src_data[106]~combout ),
	.src_data_107(\mm_interconnect_0|rsp_mux_001|src_data[107]~combout ),
	.src_data_108(\mm_interconnect_0|rsp_mux_001|src_data[108]~combout ),
	.src_payload34(\mm_interconnect_0|rsp_mux_001|src_payload~75_combout ),
	.src_data_110(\mm_interconnect_0|rsp_mux_001|src_data[110]~combout ),
	.src_data_111(\mm_interconnect_0|rsp_mux_001|src_data[111]~combout ),
	.src_data_112(\mm_interconnect_0|rsp_mux_001|src_data[112]~combout ),
	.src_payload35(\mm_interconnect_0|rsp_mux_001|src_payload~76_combout ),
	.src_data_114(\mm_interconnect_0|rsp_mux_001|src_data[114]~combout ),
	.src_data_115(\mm_interconnect_0|rsp_mux_001|src_data[115]~combout ),
	.src_payload36(\mm_interconnect_0|rsp_mux_001|src_payload~77_combout ),
	.src_data_117(\mm_interconnect_0|rsp_mux_001|src_data[117]~combout ),
	.src_payload37(\mm_interconnect_0|rsp_mux_001|src_payload~78_combout ),
	.src_data_119(\mm_interconnect_0|rsp_mux_001|src_data[119]~combout ),
	.src_payload38(\mm_interconnect_0|rsp_mux_001|src_payload~79_combout ),
	.src_data_121(\mm_interconnect_0|rsp_mux_001|src_data[121]~combout ),
	.src_data_122(\mm_interconnect_0|rsp_mux_001|src_data[122]~combout ),
	.src_data_123(\mm_interconnect_0|rsp_mux_001|src_data[123]~combout ),
	.src_data_124(\mm_interconnect_0|rsp_mux_001|src_data[124]~combout ),
	.src_payload39(\mm_interconnect_0|rsp_mux_001|src_payload~80_combout ),
	.src_data_126(\mm_interconnect_0|rsp_mux_001|src_data[126]~combout ),
	.src_data_127(\mm_interconnect_0|rsp_mux_001|src_data[127]~combout ),
	.src_data_2091(\mm_interconnect_0|rsp_mux_001|src_data[209]~combout ),
	.src_data_2101(\mm_interconnect_0|rsp_mux_001|src_data[210]~combout ),
	.src_data_2111(\mm_interconnect_0|rsp_mux_001|src_data[211]~combout ),
	.src_data_2121(\mm_interconnect_0|rsp_mux_001|src_data[212]~combout ),
	.src_data_2131(\mm_interconnect_0|rsp_mux_001|src_data[213]~combout ),
	.src_data_2141(\mm_interconnect_0|rsp_mux_001|src_data[214]~combout ),
	.src_data_2151(\mm_interconnect_0|rsp_mux_001|src_data[215]~combout ),
	.src_data_2161(\mm_interconnect_0|rsp_mux_001|src_data[216]~combout ),
	.src_data_2171(\mm_interconnect_0|rsp_mux_001|src_data[217]~combout ),
	.src_data_2181(\mm_interconnect_0|rsp_mux_001|src_data[218]~combout ),
	.src_data_2191(\mm_interconnect_0|rsp_mux_001|src_data[219]~combout ),
	.src_data_2201(\mm_interconnect_0|rsp_mux_001|src_data[220]~combout ),
	.m0_write(\mm_interconnect_0|fifo_hps_to_fpga_in_agent|m0_write~0_combout ),
	.in_data_reg_0(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.in_data_reg_1(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_2(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_3(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_4(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_5(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_6(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_7(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_8(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_9(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_10(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_11(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_12(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_13(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_14(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_15(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_16(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_17(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_18(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_19(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_20(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_21(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_22(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_23(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_24(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.in_data_reg_25(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_26(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_27(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_28(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_29(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_30(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_31(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.m0_write1(\mm_interconnect_0|onchip_sram_s2_agent|m0_write~0_combout ),
	.in_data_reg_01(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.in_data_reg_110(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_210(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_32(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_41(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_51(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_61(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_71(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_81(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_91(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_101(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_111(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_121(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_131(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_141(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_151(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_161(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_171(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_181(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_191(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_201(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_211(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_221(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_231(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_241(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.in_data_reg_251(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_261(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_271(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_281(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_291(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_301(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_311(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.r_sync_rst(\rst_controller_001|r_sync_rst~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.wrfull3(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~4_combout ),
	.wrfull4(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~5_combout ));

Computer_System_Computer_System_fifo_HPS_to_FPGA fifo_hps_to_fpga(
	.q_b_0(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[0] ),
	.q_b_1(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[1] ),
	.q_b_2(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[2] ),
	.q_b_3(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[3] ),
	.q_b_4(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[4] ),
	.q_b_5(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[5] ),
	.q_b_6(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[6] ),
	.q_b_7(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[7] ),
	.q_b_8(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[8] ),
	.q_b_9(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[9] ),
	.q_b_10(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[10] ),
	.q_b_11(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[11] ),
	.q_b_12(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[12] ),
	.q_b_13(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[13] ),
	.q_b_14(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[14] ),
	.q_b_15(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[15] ),
	.q_b_16(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[16] ),
	.q_b_17(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[17] ),
	.q_b_18(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[18] ),
	.q_b_19(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[19] ),
	.q_b_20(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[20] ),
	.q_b_21(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[21] ),
	.q_b_22(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[22] ),
	.q_b_23(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[23] ),
	.q_b_24(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[24] ),
	.q_b_25(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[25] ),
	.q_b_26(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[26] ),
	.q_b_27(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[27] ),
	.q_b_28(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[28] ),
	.q_b_29(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[29] ),
	.q_b_30(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[30] ),
	.q_b_31(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[31] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.op_2(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|op_2~13_sumout ),
	.op_21(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|op_2~25_sumout ),
	.op_22(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|op_2~29_sumout ),
	.aneb_result_wire_0(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~combout ),
	.rdclk_control_slave_readdata_0(\fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[0]~q ),
	.rdclk_control_slave_readdata_1(\fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[1]~q ),
	.rdclk_control_slave_readdata_2(\fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[2]~q ),
	.rdclk_control_slave_readdata_3(\fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[3]~q ),
	.rdclk_control_slave_readdata_4(\fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[4]~q ),
	.rdclk_control_slave_readdata_5(\fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[5]~q ),
	.rdclk_control_slave_readdata_6(\fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[6]~q ),
	.rdclk_control_slave_readdata_7(\fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[7]~q ),
	.wait_latency_counter_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_1(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_translator|wait_latency_counter[1]~q ),
	.avalonmm_write_slave_waitrequest(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~0_combout ),
	.wrfull(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~1_combout ),
	.wrfull1(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~2_combout ),
	.m0_write(\mm_interconnect_0|fifo_hps_to_fpga_in_agent|m0_write~0_combout ),
	.in_data_reg_0(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.in_data_reg_1(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_2(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_3(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_4(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_5(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_6(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_7(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_8(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_9(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_10(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_11(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_12(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_13(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_14(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_15(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_16(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_17(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_18(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_19(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_20(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_21(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_22(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_23(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_24(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.in_data_reg_25(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_26(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_27(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_28(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_29(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_30(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_31(\mm_interconnect_0|fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.r_sync_rst1(\rst_controller_001|r_sync_rst~q ),
	.m0_write1(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent|m0_write~combout ),
	.m0_read(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent|m0_read~0_combout ),
	.wrclk_control_slave_readdata_0(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[0]~q ),
	.wrclk_control_slave_readdata_1(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[1]~q ),
	.wrclk_control_slave_readdata_2(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[2]~q ),
	.wrclk_control_slave_readdata_3(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[3]~q ),
	.wrclk_control_slave_readdata_4(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[4]~q ),
	.wrclk_control_slave_readdata_5(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[5]~q ),
	.wrclk_control_slave_readdata_6(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[6]~q ),
	.wrclk_control_slave_readdata_7(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[7]~q ),
	.wrfull2(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~4_combout ),
	.wrfull3(\fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|wrfull~5_combout ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_4(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.in_data_reg_01(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.in_data_reg_210(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_110(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_141(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_81(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_131(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_121(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_111(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_101(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_91(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_191(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_181(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_171(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_161(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_151(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_261(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_211(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_201(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_311(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.in_data_reg_301(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_291(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_281(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_271(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_251(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_241(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.in_data_reg_231(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_221(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_71(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_61(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_51(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_41(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_32(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.fifo_hps_to_fpga_out_read(\fifo_hps_to_fpga_out_read~input_o ),
	.clock_bridge_0_in_clk_clk(\clock_bridge_0_in_clk_clk~input_o ),
	.fifo_hps_to_fpga_out_csr_address_2(\fifo_hps_to_fpga_out_csr_address[2]~input_o ),
	.fifo_hps_to_fpga_out_csr_address_0(\fifo_hps_to_fpga_out_csr_address[0]~input_o ),
	.fifo_hps_to_fpga_out_csr_address_1(\fifo_hps_to_fpga_out_csr_address[1]~input_o ),
	.fifo_hps_to_fpga_out_csr_read(\fifo_hps_to_fpga_out_csr_read~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_0(\fifo_hps_to_fpga_out_csr_writedata[0]~input_o ),
	.fifo_hps_to_fpga_out_csr_write(\fifo_hps_to_fpga_out_csr_write~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_7(\fifo_hps_to_fpga_out_csr_writedata[7]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_1(\fifo_hps_to_fpga_out_csr_writedata[1]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_13(\fifo_hps_to_fpga_out_csr_writedata[13]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_19(\fifo_hps_to_fpga_out_csr_writedata[19]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_26(\fifo_hps_to_fpga_out_csr_writedata[26]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_27(\fifo_hps_to_fpga_out_csr_writedata[27]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_28(\fifo_hps_to_fpga_out_csr_writedata[28]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_29(\fifo_hps_to_fpga_out_csr_writedata[29]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_30(\fifo_hps_to_fpga_out_csr_writedata[30]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_31(\fifo_hps_to_fpga_out_csr_writedata[31]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_20(\fifo_hps_to_fpga_out_csr_writedata[20]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_21(\fifo_hps_to_fpga_out_csr_writedata[21]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_22(\fifo_hps_to_fpga_out_csr_writedata[22]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_23(\fifo_hps_to_fpga_out_csr_writedata[23]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_24(\fifo_hps_to_fpga_out_csr_writedata[24]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_25(\fifo_hps_to_fpga_out_csr_writedata[25]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_8(\fifo_hps_to_fpga_out_csr_writedata[8]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_9(\fifo_hps_to_fpga_out_csr_writedata[9]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_10(\fifo_hps_to_fpga_out_csr_writedata[10]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_11(\fifo_hps_to_fpga_out_csr_writedata[11]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_12(\fifo_hps_to_fpga_out_csr_writedata[12]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_14(\fifo_hps_to_fpga_out_csr_writedata[14]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_15(\fifo_hps_to_fpga_out_csr_writedata[15]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_16(\fifo_hps_to_fpga_out_csr_writedata[16]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_17(\fifo_hps_to_fpga_out_csr_writedata[17]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_18(\fifo_hps_to_fpga_out_csr_writedata[18]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_2(\fifo_hps_to_fpga_out_csr_writedata[2]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_3(\fifo_hps_to_fpga_out_csr_writedata[3]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_4(\fifo_hps_to_fpga_out_csr_writedata[4]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_5(\fifo_hps_to_fpga_out_csr_writedata[5]~input_o ),
	.fifo_hps_to_fpga_out_csr_writedata_6(\fifo_hps_to_fpga_out_csr_writedata[6]~input_o ));

Computer_System_Computer_System_System_PLL system_pll(
	.outclk_wire_1(\system_pll|sys_pll|altera_pll_i|outclk_wire[1] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.locked_wire_0(\system_pll|sys_pll|altera_pll_i|locked_wire[0] ),
	.system_pll_ref_clk_clk(\system_pll_ref_clk_clk~input_o ),
	.system_pll_ref_reset_reset(\system_pll_ref_reset_reset~input_o ));

Computer_System_Computer_System_Onchip_SRAM onchip_sram(
	.q_a_0(\onchip_sram|the_altsyncram|auto_generated|q_a[0] ),
	.q_b_0(\onchip_sram|the_altsyncram|auto_generated|q_b[0] ),
	.q_a_1(\onchip_sram|the_altsyncram|auto_generated|q_a[1] ),
	.q_b_1(\onchip_sram|the_altsyncram|auto_generated|q_b[1] ),
	.q_a_2(\onchip_sram|the_altsyncram|auto_generated|q_a[2] ),
	.q_b_2(\onchip_sram|the_altsyncram|auto_generated|q_b[2] ),
	.q_a_3(\onchip_sram|the_altsyncram|auto_generated|q_a[3] ),
	.q_b_3(\onchip_sram|the_altsyncram|auto_generated|q_b[3] ),
	.q_a_4(\onchip_sram|the_altsyncram|auto_generated|q_a[4] ),
	.q_b_4(\onchip_sram|the_altsyncram|auto_generated|q_b[4] ),
	.q_a_5(\onchip_sram|the_altsyncram|auto_generated|q_a[5] ),
	.q_b_5(\onchip_sram|the_altsyncram|auto_generated|q_b[5] ),
	.q_a_6(\onchip_sram|the_altsyncram|auto_generated|q_a[6] ),
	.q_b_6(\onchip_sram|the_altsyncram|auto_generated|q_b[6] ),
	.q_a_7(\onchip_sram|the_altsyncram|auto_generated|q_a[7] ),
	.q_b_7(\onchip_sram|the_altsyncram|auto_generated|q_b[7] ),
	.q_a_8(\onchip_sram|the_altsyncram|auto_generated|q_a[8] ),
	.q_b_8(\onchip_sram|the_altsyncram|auto_generated|q_b[8] ),
	.q_a_9(\onchip_sram|the_altsyncram|auto_generated|q_a[9] ),
	.q_b_9(\onchip_sram|the_altsyncram|auto_generated|q_b[9] ),
	.q_a_10(\onchip_sram|the_altsyncram|auto_generated|q_a[10] ),
	.q_b_10(\onchip_sram|the_altsyncram|auto_generated|q_b[10] ),
	.q_a_11(\onchip_sram|the_altsyncram|auto_generated|q_a[11] ),
	.q_b_11(\onchip_sram|the_altsyncram|auto_generated|q_b[11] ),
	.q_a_12(\onchip_sram|the_altsyncram|auto_generated|q_a[12] ),
	.q_b_12(\onchip_sram|the_altsyncram|auto_generated|q_b[12] ),
	.q_a_13(\onchip_sram|the_altsyncram|auto_generated|q_a[13] ),
	.q_b_13(\onchip_sram|the_altsyncram|auto_generated|q_b[13] ),
	.q_a_14(\onchip_sram|the_altsyncram|auto_generated|q_a[14] ),
	.q_b_14(\onchip_sram|the_altsyncram|auto_generated|q_b[14] ),
	.q_a_15(\onchip_sram|the_altsyncram|auto_generated|q_a[15] ),
	.q_b_15(\onchip_sram|the_altsyncram|auto_generated|q_b[15] ),
	.q_a_16(\onchip_sram|the_altsyncram|auto_generated|q_a[16] ),
	.q_b_16(\onchip_sram|the_altsyncram|auto_generated|q_b[16] ),
	.q_a_17(\onchip_sram|the_altsyncram|auto_generated|q_a[17] ),
	.q_b_17(\onchip_sram|the_altsyncram|auto_generated|q_b[17] ),
	.q_a_18(\onchip_sram|the_altsyncram|auto_generated|q_a[18] ),
	.q_b_18(\onchip_sram|the_altsyncram|auto_generated|q_b[18] ),
	.q_a_19(\onchip_sram|the_altsyncram|auto_generated|q_a[19] ),
	.q_b_19(\onchip_sram|the_altsyncram|auto_generated|q_b[19] ),
	.q_a_20(\onchip_sram|the_altsyncram|auto_generated|q_a[20] ),
	.q_b_20(\onchip_sram|the_altsyncram|auto_generated|q_b[20] ),
	.q_a_21(\onchip_sram|the_altsyncram|auto_generated|q_a[21] ),
	.q_b_21(\onchip_sram|the_altsyncram|auto_generated|q_b[21] ),
	.q_a_22(\onchip_sram|the_altsyncram|auto_generated|q_a[22] ),
	.q_b_22(\onchip_sram|the_altsyncram|auto_generated|q_b[22] ),
	.q_a_23(\onchip_sram|the_altsyncram|auto_generated|q_a[23] ),
	.q_b_23(\onchip_sram|the_altsyncram|auto_generated|q_b[23] ),
	.q_a_24(\onchip_sram|the_altsyncram|auto_generated|q_a[24] ),
	.q_b_24(\onchip_sram|the_altsyncram|auto_generated|q_b[24] ),
	.q_a_25(\onchip_sram|the_altsyncram|auto_generated|q_a[25] ),
	.q_b_25(\onchip_sram|the_altsyncram|auto_generated|q_b[25] ),
	.q_a_26(\onchip_sram|the_altsyncram|auto_generated|q_a[26] ),
	.q_b_26(\onchip_sram|the_altsyncram|auto_generated|q_b[26] ),
	.q_a_27(\onchip_sram|the_altsyncram|auto_generated|q_a[27] ),
	.q_b_27(\onchip_sram|the_altsyncram|auto_generated|q_b[27] ),
	.q_a_28(\onchip_sram|the_altsyncram|auto_generated|q_a[28] ),
	.q_b_28(\onchip_sram|the_altsyncram|auto_generated|q_b[28] ),
	.q_a_29(\onchip_sram|the_altsyncram|auto_generated|q_a[29] ),
	.q_b_29(\onchip_sram|the_altsyncram|auto_generated|q_b[29] ),
	.q_a_30(\onchip_sram|the_altsyncram|auto_generated|q_a[30] ),
	.q_b_30(\onchip_sram|the_altsyncram|auto_generated|q_b[30] ),
	.q_a_31(\onchip_sram|the_altsyncram|auto_generated|q_a[31] ),
	.q_b_31(\onchip_sram|the_altsyncram|auto_generated|q_b[31] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_4(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ),
	.int_nxt_addr_reg_dly_5(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[5]~q ),
	.int_nxt_addr_reg_dly_6(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[6]~q ),
	.int_nxt_addr_reg_dly_7(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[7]~q ),
	.int_nxt_addr_reg_dly_8(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[8]~q ),
	.int_nxt_addr_reg_dly_9(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[9]~q ),
	.source0_data_34(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[34]~0_combout ),
	.source0_data_32(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[32]~1_combout ),
	.source0_data_33(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[33]~2_combout ),
	.source0_data_35(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~4_combout ),
	.m0_write(\mm_interconnect_0|onchip_sram_s2_agent|m0_write~0_combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.r_early_rst1(\rst_controller_001|r_early_rst~q ),
	.in_data_reg_0(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.in_data_reg_1(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_2(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_3(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_4(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_5(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_6(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_7(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_8(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_9(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_10(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_11(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_12(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_13(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_14(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_15(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_16(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_17(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_18(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_19(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_20(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_21(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_22(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_23(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_24(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.in_data_reg_25(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_26(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_27(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_28(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_29(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_30(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_31(\mm_interconnect_0|onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.clock_bridge_0_in_clk_clk(\clock_bridge_0_in_clk_clk~input_o ),
	.onchip_sram_s1_chipselect(\onchip_sram_s1_chipselect~input_o ),
	.onchip_sram_s1_write(\onchip_sram_s1_write~input_o ),
	.onchip_sram_s1_clken(\onchip_sram_s1_clken~input_o ),
	.onchip_sram_s1_writedata_0(\onchip_sram_s1_writedata[0]~input_o ),
	.onchip_sram_s1_address_0(\onchip_sram_s1_address[0]~input_o ),
	.onchip_sram_s1_address_1(\onchip_sram_s1_address[1]~input_o ),
	.onchip_sram_s1_address_2(\onchip_sram_s1_address[2]~input_o ),
	.onchip_sram_s1_address_3(\onchip_sram_s1_address[3]~input_o ),
	.onchip_sram_s1_address_4(\onchip_sram_s1_address[4]~input_o ),
	.onchip_sram_s1_address_5(\onchip_sram_s1_address[5]~input_o ),
	.onchip_sram_s1_address_6(\onchip_sram_s1_address[6]~input_o ),
	.onchip_sram_s1_address_7(\onchip_sram_s1_address[7]~input_o ),
	.onchip_sram_s1_byteenable_0(\onchip_sram_s1_byteenable[0]~input_o ),
	.onchip_sram_s1_writedata_1(\onchip_sram_s1_writedata[1]~input_o ),
	.onchip_sram_s1_writedata_2(\onchip_sram_s1_writedata[2]~input_o ),
	.onchip_sram_s1_writedata_3(\onchip_sram_s1_writedata[3]~input_o ),
	.onchip_sram_s1_writedata_4(\onchip_sram_s1_writedata[4]~input_o ),
	.onchip_sram_s1_writedata_5(\onchip_sram_s1_writedata[5]~input_o ),
	.onchip_sram_s1_writedata_6(\onchip_sram_s1_writedata[6]~input_o ),
	.onchip_sram_s1_writedata_7(\onchip_sram_s1_writedata[7]~input_o ),
	.onchip_sram_s1_writedata_8(\onchip_sram_s1_writedata[8]~input_o ),
	.onchip_sram_s1_byteenable_1(\onchip_sram_s1_byteenable[1]~input_o ),
	.onchip_sram_s1_writedata_9(\onchip_sram_s1_writedata[9]~input_o ),
	.onchip_sram_s1_writedata_10(\onchip_sram_s1_writedata[10]~input_o ),
	.onchip_sram_s1_writedata_11(\onchip_sram_s1_writedata[11]~input_o ),
	.onchip_sram_s1_writedata_12(\onchip_sram_s1_writedata[12]~input_o ),
	.onchip_sram_s1_writedata_13(\onchip_sram_s1_writedata[13]~input_o ),
	.onchip_sram_s1_writedata_14(\onchip_sram_s1_writedata[14]~input_o ),
	.onchip_sram_s1_writedata_15(\onchip_sram_s1_writedata[15]~input_o ),
	.onchip_sram_s1_writedata_16(\onchip_sram_s1_writedata[16]~input_o ),
	.onchip_sram_s1_byteenable_2(\onchip_sram_s1_byteenable[2]~input_o ),
	.onchip_sram_s1_writedata_17(\onchip_sram_s1_writedata[17]~input_o ),
	.onchip_sram_s1_writedata_18(\onchip_sram_s1_writedata[18]~input_o ),
	.onchip_sram_s1_writedata_19(\onchip_sram_s1_writedata[19]~input_o ),
	.onchip_sram_s1_writedata_20(\onchip_sram_s1_writedata[20]~input_o ),
	.onchip_sram_s1_writedata_21(\onchip_sram_s1_writedata[21]~input_o ),
	.onchip_sram_s1_writedata_22(\onchip_sram_s1_writedata[22]~input_o ),
	.onchip_sram_s1_writedata_23(\onchip_sram_s1_writedata[23]~input_o ),
	.onchip_sram_s1_writedata_24(\onchip_sram_s1_writedata[24]~input_o ),
	.onchip_sram_s1_byteenable_3(\onchip_sram_s1_byteenable[3]~input_o ),
	.onchip_sram_s1_writedata_25(\onchip_sram_s1_writedata[25]~input_o ),
	.onchip_sram_s1_writedata_26(\onchip_sram_s1_writedata[26]~input_o ),
	.onchip_sram_s1_writedata_27(\onchip_sram_s1_writedata[27]~input_o ),
	.onchip_sram_s1_writedata_28(\onchip_sram_s1_writedata[28]~input_o ),
	.onchip_sram_s1_writedata_29(\onchip_sram_s1_writedata[29]~input_o ),
	.onchip_sram_s1_writedata_30(\onchip_sram_s1_writedata[30]~input_o ),
	.onchip_sram_s1_writedata_31(\onchip_sram_s1_writedata[31]~input_o ));

Computer_System_Computer_System_ARM_A9_HPS arm_a9_hps(
	.h2f_rst_n_0(\arm_a9_hps|fpga_interfaces|h2f_rst_n[0] ),
	.h2f_lw_ARVALID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARVALID[0] ),
	.h2f_lw_AWVALID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWVALID[0] ),
	.h2f_lw_BREADY_0(\arm_a9_hps|fpga_interfaces|h2f_lw_BREADY[0] ),
	.h2f_lw_RREADY_0(\arm_a9_hps|fpga_interfaces|h2f_lw_RREADY[0] ),
	.h2f_lw_WLAST_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WLAST[0] ),
	.h2f_lw_WVALID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WVALID[0] ),
	.h2f_lw_ARADDR_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[0] ),
	.h2f_lw_ARADDR_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[1] ),
	.h2f_lw_ARADDR_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[2] ),
	.h2f_lw_ARADDR_3(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[3] ),
	.h2f_lw_ARADDR_4(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[4] ),
	.h2f_lw_ARBURST_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARBURST[0] ),
	.h2f_lw_ARBURST_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARBURST[1] ),
	.h2f_lw_ARID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[0] ),
	.h2f_lw_ARID_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[1] ),
	.h2f_lw_ARID_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[2] ),
	.h2f_lw_ARID_3(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[3] ),
	.h2f_lw_ARID_4(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[4] ),
	.h2f_lw_ARID_5(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[5] ),
	.h2f_lw_ARID_6(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[6] ),
	.h2f_lw_ARID_7(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[7] ),
	.h2f_lw_ARID_8(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[8] ),
	.h2f_lw_ARID_9(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[9] ),
	.h2f_lw_ARID_10(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[10] ),
	.h2f_lw_ARID_11(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[11] ),
	.h2f_lw_ARLEN_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[0] ),
	.h2f_lw_ARLEN_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[1] ),
	.h2f_lw_ARLEN_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[2] ),
	.h2f_lw_ARLEN_3(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[3] ),
	.h2f_lw_ARSIZE_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[0] ),
	.h2f_lw_ARSIZE_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[1] ),
	.h2f_lw_ARSIZE_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[2] ),
	.h2f_lw_AWADDR_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[0] ),
	.h2f_lw_AWADDR_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[1] ),
	.h2f_lw_AWADDR_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[2] ),
	.h2f_lw_AWADDR_3(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[3] ),
	.h2f_lw_AWADDR_4(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[4] ),
	.h2f_lw_AWBURST_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWBURST[0] ),
	.h2f_lw_AWBURST_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWBURST[1] ),
	.h2f_lw_AWID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[0] ),
	.h2f_lw_AWID_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[1] ),
	.h2f_lw_AWID_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[2] ),
	.h2f_lw_AWID_3(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[3] ),
	.h2f_lw_AWID_4(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[4] ),
	.h2f_lw_AWID_5(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[5] ),
	.h2f_lw_AWID_6(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[6] ),
	.h2f_lw_AWID_7(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[7] ),
	.h2f_lw_AWID_8(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[8] ),
	.h2f_lw_AWID_9(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[9] ),
	.h2f_lw_AWID_10(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[10] ),
	.h2f_lw_AWID_11(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[11] ),
	.h2f_lw_AWLEN_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[0] ),
	.h2f_lw_AWLEN_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[1] ),
	.h2f_lw_AWLEN_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[2] ),
	.h2f_lw_AWLEN_3(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[3] ),
	.h2f_lw_AWSIZE_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[0] ),
	.h2f_lw_AWSIZE_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[1] ),
	.h2f_lw_AWSIZE_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[2] ),
	.h2f_lw_WDATA_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[0] ),
	.h2f_lw_WDATA_1(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[1] ),
	.h2f_lw_WDATA_2(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[2] ),
	.h2f_lw_WDATA_3(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[3] ),
	.h2f_lw_WDATA_4(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[4] ),
	.h2f_lw_WDATA_5(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[5] ),
	.h2f_lw_WDATA_6(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[6] ),
	.h2f_lw_WDATA_7(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[7] ),
	.h2f_lw_WDATA_8(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[8] ),
	.h2f_lw_WDATA_9(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[9] ),
	.h2f_lw_WDATA_10(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[10] ),
	.h2f_lw_WDATA_11(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[11] ),
	.h2f_lw_WDATA_12(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[12] ),
	.h2f_lw_WDATA_13(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[13] ),
	.h2f_lw_WDATA_14(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[14] ),
	.h2f_lw_WDATA_15(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[15] ),
	.h2f_lw_WDATA_16(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[16] ),
	.h2f_lw_WDATA_17(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[17] ),
	.h2f_lw_WDATA_18(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[18] ),
	.h2f_lw_WDATA_19(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[19] ),
	.h2f_lw_WDATA_20(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[20] ),
	.h2f_lw_WDATA_21(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[21] ),
	.h2f_lw_WDATA_22(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[22] ),
	.h2f_lw_WDATA_23(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[23] ),
	.h2f_lw_WDATA_24(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[24] ),
	.h2f_lw_WDATA_25(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[25] ),
	.h2f_lw_WDATA_26(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[26] ),
	.h2f_lw_WDATA_27(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[27] ),
	.h2f_lw_WDATA_28(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[28] ),
	.h2f_lw_WDATA_29(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[29] ),
	.h2f_lw_WDATA_30(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[30] ),
	.h2f_lw_WDATA_31(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[31] ),
	.h2f_lw_WSTRB_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[0] ),
	.h2f_lw_WSTRB_1(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[1] ),
	.h2f_lw_WSTRB_2(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[2] ),
	.h2f_lw_WSTRB_3(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[3] ),
	.h2f_ARVALID_0(\arm_a9_hps|fpga_interfaces|h2f_ARVALID[0] ),
	.h2f_AWVALID_0(\arm_a9_hps|fpga_interfaces|h2f_AWVALID[0] ),
	.h2f_BREADY_0(\arm_a9_hps|fpga_interfaces|h2f_BREADY[0] ),
	.h2f_RREADY_0(\arm_a9_hps|fpga_interfaces|h2f_RREADY[0] ),
	.h2f_WLAST_0(\arm_a9_hps|fpga_interfaces|h2f_WLAST[0] ),
	.h2f_WVALID_0(\arm_a9_hps|fpga_interfaces|h2f_WVALID[0] ),
	.h2f_ARADDR_0(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[0] ),
	.h2f_ARADDR_1(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[1] ),
	.h2f_ARADDR_2(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[2] ),
	.h2f_ARADDR_3(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[3] ),
	.h2f_ARADDR_4(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[4] ),
	.h2f_ARADDR_5(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[5] ),
	.h2f_ARADDR_6(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[6] ),
	.h2f_ARADDR_7(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[7] ),
	.h2f_ARADDR_8(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[8] ),
	.h2f_ARADDR_9(\arm_a9_hps|fpga_interfaces|h2f_ARADDR[9] ),
	.h2f_ARBURST_0(\arm_a9_hps|fpga_interfaces|h2f_ARBURST[0] ),
	.h2f_ARBURST_1(\arm_a9_hps|fpga_interfaces|h2f_ARBURST[1] ),
	.h2f_ARID_0(\arm_a9_hps|fpga_interfaces|h2f_ARID[0] ),
	.h2f_ARID_1(\arm_a9_hps|fpga_interfaces|h2f_ARID[1] ),
	.h2f_ARID_2(\arm_a9_hps|fpga_interfaces|h2f_ARID[2] ),
	.h2f_ARID_3(\arm_a9_hps|fpga_interfaces|h2f_ARID[3] ),
	.h2f_ARID_4(\arm_a9_hps|fpga_interfaces|h2f_ARID[4] ),
	.h2f_ARID_5(\arm_a9_hps|fpga_interfaces|h2f_ARID[5] ),
	.h2f_ARID_6(\arm_a9_hps|fpga_interfaces|h2f_ARID[6] ),
	.h2f_ARID_7(\arm_a9_hps|fpga_interfaces|h2f_ARID[7] ),
	.h2f_ARID_8(\arm_a9_hps|fpga_interfaces|h2f_ARID[8] ),
	.h2f_ARID_9(\arm_a9_hps|fpga_interfaces|h2f_ARID[9] ),
	.h2f_ARID_10(\arm_a9_hps|fpga_interfaces|h2f_ARID[10] ),
	.h2f_ARID_11(\arm_a9_hps|fpga_interfaces|h2f_ARID[11] ),
	.h2f_ARLEN_0(\arm_a9_hps|fpga_interfaces|h2f_ARLEN[0] ),
	.h2f_ARLEN_1(\arm_a9_hps|fpga_interfaces|h2f_ARLEN[1] ),
	.h2f_ARLEN_2(\arm_a9_hps|fpga_interfaces|h2f_ARLEN[2] ),
	.h2f_ARLEN_3(\arm_a9_hps|fpga_interfaces|h2f_ARLEN[3] ),
	.h2f_ARSIZE_0(\arm_a9_hps|fpga_interfaces|h2f_ARSIZE[0] ),
	.h2f_ARSIZE_1(\arm_a9_hps|fpga_interfaces|h2f_ARSIZE[1] ),
	.h2f_ARSIZE_2(\arm_a9_hps|fpga_interfaces|h2f_ARSIZE[2] ),
	.h2f_AWADDR_0(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[0] ),
	.h2f_AWADDR_1(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[1] ),
	.h2f_AWADDR_2(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[2] ),
	.h2f_AWADDR_3(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[3] ),
	.h2f_AWADDR_4(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[4] ),
	.h2f_AWADDR_5(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[5] ),
	.h2f_AWADDR_6(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[6] ),
	.h2f_AWADDR_7(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[7] ),
	.h2f_AWADDR_8(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[8] ),
	.h2f_AWADDR_9(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[9] ),
	.h2f_AWADDR_10(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[10] ),
	.h2f_AWADDR_11(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[11] ),
	.h2f_AWADDR_12(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[12] ),
	.h2f_AWADDR_13(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[13] ),
	.h2f_AWADDR_14(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[14] ),
	.h2f_AWADDR_15(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[15] ),
	.h2f_AWADDR_16(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[16] ),
	.h2f_AWADDR_17(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[17] ),
	.h2f_AWADDR_18(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[18] ),
	.h2f_AWADDR_19(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[19] ),
	.h2f_AWADDR_20(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[20] ),
	.h2f_AWADDR_21(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[21] ),
	.h2f_AWADDR_22(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[22] ),
	.h2f_AWADDR_23(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[23] ),
	.h2f_AWADDR_24(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[24] ),
	.h2f_AWADDR_25(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[25] ),
	.h2f_AWADDR_26(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[26] ),
	.h2f_AWADDR_27(\arm_a9_hps|fpga_interfaces|h2f_AWADDR[27] ),
	.h2f_AWBURST_0(\arm_a9_hps|fpga_interfaces|h2f_AWBURST[0] ),
	.h2f_AWBURST_1(\arm_a9_hps|fpga_interfaces|h2f_AWBURST[1] ),
	.h2f_AWID_0(\arm_a9_hps|fpga_interfaces|h2f_AWID[0] ),
	.h2f_AWID_1(\arm_a9_hps|fpga_interfaces|h2f_AWID[1] ),
	.h2f_AWID_2(\arm_a9_hps|fpga_interfaces|h2f_AWID[2] ),
	.h2f_AWID_3(\arm_a9_hps|fpga_interfaces|h2f_AWID[3] ),
	.h2f_AWID_4(\arm_a9_hps|fpga_interfaces|h2f_AWID[4] ),
	.h2f_AWID_5(\arm_a9_hps|fpga_interfaces|h2f_AWID[5] ),
	.h2f_AWID_6(\arm_a9_hps|fpga_interfaces|h2f_AWID[6] ),
	.h2f_AWID_7(\arm_a9_hps|fpga_interfaces|h2f_AWID[7] ),
	.h2f_AWID_8(\arm_a9_hps|fpga_interfaces|h2f_AWID[8] ),
	.h2f_AWID_9(\arm_a9_hps|fpga_interfaces|h2f_AWID[9] ),
	.h2f_AWID_10(\arm_a9_hps|fpga_interfaces|h2f_AWID[10] ),
	.h2f_AWID_11(\arm_a9_hps|fpga_interfaces|h2f_AWID[11] ),
	.h2f_AWLEN_0(\arm_a9_hps|fpga_interfaces|h2f_AWLEN[0] ),
	.h2f_AWLEN_1(\arm_a9_hps|fpga_interfaces|h2f_AWLEN[1] ),
	.h2f_AWLEN_2(\arm_a9_hps|fpga_interfaces|h2f_AWLEN[2] ),
	.h2f_AWLEN_3(\arm_a9_hps|fpga_interfaces|h2f_AWLEN[3] ),
	.h2f_AWSIZE_0(\arm_a9_hps|fpga_interfaces|h2f_AWSIZE[0] ),
	.h2f_AWSIZE_1(\arm_a9_hps|fpga_interfaces|h2f_AWSIZE[1] ),
	.h2f_AWSIZE_2(\arm_a9_hps|fpga_interfaces|h2f_AWSIZE[2] ),
	.h2f_WDATA_0(\arm_a9_hps|fpga_interfaces|h2f_WDATA[0] ),
	.h2f_WDATA_1(\arm_a9_hps|fpga_interfaces|h2f_WDATA[1] ),
	.h2f_WDATA_2(\arm_a9_hps|fpga_interfaces|h2f_WDATA[2] ),
	.h2f_WDATA_3(\arm_a9_hps|fpga_interfaces|h2f_WDATA[3] ),
	.h2f_WDATA_4(\arm_a9_hps|fpga_interfaces|h2f_WDATA[4] ),
	.h2f_WDATA_5(\arm_a9_hps|fpga_interfaces|h2f_WDATA[5] ),
	.h2f_WDATA_6(\arm_a9_hps|fpga_interfaces|h2f_WDATA[6] ),
	.h2f_WDATA_7(\arm_a9_hps|fpga_interfaces|h2f_WDATA[7] ),
	.h2f_WDATA_8(\arm_a9_hps|fpga_interfaces|h2f_WDATA[8] ),
	.h2f_WDATA_9(\arm_a9_hps|fpga_interfaces|h2f_WDATA[9] ),
	.h2f_WDATA_10(\arm_a9_hps|fpga_interfaces|h2f_WDATA[10] ),
	.h2f_WDATA_11(\arm_a9_hps|fpga_interfaces|h2f_WDATA[11] ),
	.h2f_WDATA_12(\arm_a9_hps|fpga_interfaces|h2f_WDATA[12] ),
	.h2f_WDATA_13(\arm_a9_hps|fpga_interfaces|h2f_WDATA[13] ),
	.h2f_WDATA_14(\arm_a9_hps|fpga_interfaces|h2f_WDATA[14] ),
	.h2f_WDATA_15(\arm_a9_hps|fpga_interfaces|h2f_WDATA[15] ),
	.h2f_WDATA_16(\arm_a9_hps|fpga_interfaces|h2f_WDATA[16] ),
	.h2f_WDATA_17(\arm_a9_hps|fpga_interfaces|h2f_WDATA[17] ),
	.h2f_WDATA_18(\arm_a9_hps|fpga_interfaces|h2f_WDATA[18] ),
	.h2f_WDATA_19(\arm_a9_hps|fpga_interfaces|h2f_WDATA[19] ),
	.h2f_WDATA_20(\arm_a9_hps|fpga_interfaces|h2f_WDATA[20] ),
	.h2f_WDATA_21(\arm_a9_hps|fpga_interfaces|h2f_WDATA[21] ),
	.h2f_WDATA_22(\arm_a9_hps|fpga_interfaces|h2f_WDATA[22] ),
	.h2f_WDATA_23(\arm_a9_hps|fpga_interfaces|h2f_WDATA[23] ),
	.h2f_WDATA_24(\arm_a9_hps|fpga_interfaces|h2f_WDATA[24] ),
	.h2f_WDATA_25(\arm_a9_hps|fpga_interfaces|h2f_WDATA[25] ),
	.h2f_WDATA_26(\arm_a9_hps|fpga_interfaces|h2f_WDATA[26] ),
	.h2f_WDATA_27(\arm_a9_hps|fpga_interfaces|h2f_WDATA[27] ),
	.h2f_WDATA_28(\arm_a9_hps|fpga_interfaces|h2f_WDATA[28] ),
	.h2f_WDATA_29(\arm_a9_hps|fpga_interfaces|h2f_WDATA[29] ),
	.h2f_WDATA_30(\arm_a9_hps|fpga_interfaces|h2f_WDATA[30] ),
	.h2f_WDATA_31(\arm_a9_hps|fpga_interfaces|h2f_WDATA[31] ),
	.h2f_WDATA_32(\arm_a9_hps|fpga_interfaces|h2f_WDATA[32] ),
	.h2f_WDATA_33(\arm_a9_hps|fpga_interfaces|h2f_WDATA[33] ),
	.h2f_WDATA_34(\arm_a9_hps|fpga_interfaces|h2f_WDATA[34] ),
	.h2f_WDATA_35(\arm_a9_hps|fpga_interfaces|h2f_WDATA[35] ),
	.h2f_WDATA_36(\arm_a9_hps|fpga_interfaces|h2f_WDATA[36] ),
	.h2f_WDATA_37(\arm_a9_hps|fpga_interfaces|h2f_WDATA[37] ),
	.h2f_WDATA_38(\arm_a9_hps|fpga_interfaces|h2f_WDATA[38] ),
	.h2f_WDATA_39(\arm_a9_hps|fpga_interfaces|h2f_WDATA[39] ),
	.h2f_WDATA_40(\arm_a9_hps|fpga_interfaces|h2f_WDATA[40] ),
	.h2f_WDATA_41(\arm_a9_hps|fpga_interfaces|h2f_WDATA[41] ),
	.h2f_WDATA_42(\arm_a9_hps|fpga_interfaces|h2f_WDATA[42] ),
	.h2f_WDATA_43(\arm_a9_hps|fpga_interfaces|h2f_WDATA[43] ),
	.h2f_WDATA_44(\arm_a9_hps|fpga_interfaces|h2f_WDATA[44] ),
	.h2f_WDATA_45(\arm_a9_hps|fpga_interfaces|h2f_WDATA[45] ),
	.h2f_WDATA_46(\arm_a9_hps|fpga_interfaces|h2f_WDATA[46] ),
	.h2f_WDATA_47(\arm_a9_hps|fpga_interfaces|h2f_WDATA[47] ),
	.h2f_WDATA_48(\arm_a9_hps|fpga_interfaces|h2f_WDATA[48] ),
	.h2f_WDATA_49(\arm_a9_hps|fpga_interfaces|h2f_WDATA[49] ),
	.h2f_WDATA_50(\arm_a9_hps|fpga_interfaces|h2f_WDATA[50] ),
	.h2f_WDATA_51(\arm_a9_hps|fpga_interfaces|h2f_WDATA[51] ),
	.h2f_WDATA_52(\arm_a9_hps|fpga_interfaces|h2f_WDATA[52] ),
	.h2f_WDATA_53(\arm_a9_hps|fpga_interfaces|h2f_WDATA[53] ),
	.h2f_WDATA_54(\arm_a9_hps|fpga_interfaces|h2f_WDATA[54] ),
	.h2f_WDATA_55(\arm_a9_hps|fpga_interfaces|h2f_WDATA[55] ),
	.h2f_WDATA_56(\arm_a9_hps|fpga_interfaces|h2f_WDATA[56] ),
	.h2f_WDATA_57(\arm_a9_hps|fpga_interfaces|h2f_WDATA[57] ),
	.h2f_WDATA_58(\arm_a9_hps|fpga_interfaces|h2f_WDATA[58] ),
	.h2f_WDATA_59(\arm_a9_hps|fpga_interfaces|h2f_WDATA[59] ),
	.h2f_WDATA_60(\arm_a9_hps|fpga_interfaces|h2f_WDATA[60] ),
	.h2f_WDATA_61(\arm_a9_hps|fpga_interfaces|h2f_WDATA[61] ),
	.h2f_WDATA_62(\arm_a9_hps|fpga_interfaces|h2f_WDATA[62] ),
	.h2f_WDATA_63(\arm_a9_hps|fpga_interfaces|h2f_WDATA[63] ),
	.h2f_WDATA_64(\arm_a9_hps|fpga_interfaces|h2f_WDATA[64] ),
	.h2f_WDATA_65(\arm_a9_hps|fpga_interfaces|h2f_WDATA[65] ),
	.h2f_WDATA_66(\arm_a9_hps|fpga_interfaces|h2f_WDATA[66] ),
	.h2f_WDATA_67(\arm_a9_hps|fpga_interfaces|h2f_WDATA[67] ),
	.h2f_WDATA_68(\arm_a9_hps|fpga_interfaces|h2f_WDATA[68] ),
	.h2f_WDATA_69(\arm_a9_hps|fpga_interfaces|h2f_WDATA[69] ),
	.h2f_WDATA_70(\arm_a9_hps|fpga_interfaces|h2f_WDATA[70] ),
	.h2f_WDATA_71(\arm_a9_hps|fpga_interfaces|h2f_WDATA[71] ),
	.h2f_WDATA_72(\arm_a9_hps|fpga_interfaces|h2f_WDATA[72] ),
	.h2f_WDATA_73(\arm_a9_hps|fpga_interfaces|h2f_WDATA[73] ),
	.h2f_WDATA_74(\arm_a9_hps|fpga_interfaces|h2f_WDATA[74] ),
	.h2f_WDATA_75(\arm_a9_hps|fpga_interfaces|h2f_WDATA[75] ),
	.h2f_WDATA_76(\arm_a9_hps|fpga_interfaces|h2f_WDATA[76] ),
	.h2f_WDATA_77(\arm_a9_hps|fpga_interfaces|h2f_WDATA[77] ),
	.h2f_WDATA_78(\arm_a9_hps|fpga_interfaces|h2f_WDATA[78] ),
	.h2f_WDATA_79(\arm_a9_hps|fpga_interfaces|h2f_WDATA[79] ),
	.h2f_WDATA_80(\arm_a9_hps|fpga_interfaces|h2f_WDATA[80] ),
	.h2f_WDATA_81(\arm_a9_hps|fpga_interfaces|h2f_WDATA[81] ),
	.h2f_WDATA_82(\arm_a9_hps|fpga_interfaces|h2f_WDATA[82] ),
	.h2f_WDATA_83(\arm_a9_hps|fpga_interfaces|h2f_WDATA[83] ),
	.h2f_WDATA_84(\arm_a9_hps|fpga_interfaces|h2f_WDATA[84] ),
	.h2f_WDATA_85(\arm_a9_hps|fpga_interfaces|h2f_WDATA[85] ),
	.h2f_WDATA_86(\arm_a9_hps|fpga_interfaces|h2f_WDATA[86] ),
	.h2f_WDATA_87(\arm_a9_hps|fpga_interfaces|h2f_WDATA[87] ),
	.h2f_WDATA_88(\arm_a9_hps|fpga_interfaces|h2f_WDATA[88] ),
	.h2f_WDATA_89(\arm_a9_hps|fpga_interfaces|h2f_WDATA[89] ),
	.h2f_WDATA_90(\arm_a9_hps|fpga_interfaces|h2f_WDATA[90] ),
	.h2f_WDATA_91(\arm_a9_hps|fpga_interfaces|h2f_WDATA[91] ),
	.h2f_WDATA_92(\arm_a9_hps|fpga_interfaces|h2f_WDATA[92] ),
	.h2f_WDATA_93(\arm_a9_hps|fpga_interfaces|h2f_WDATA[93] ),
	.h2f_WDATA_94(\arm_a9_hps|fpga_interfaces|h2f_WDATA[94] ),
	.h2f_WDATA_95(\arm_a9_hps|fpga_interfaces|h2f_WDATA[95] ),
	.h2f_WDATA_96(\arm_a9_hps|fpga_interfaces|h2f_WDATA[96] ),
	.h2f_WDATA_97(\arm_a9_hps|fpga_interfaces|h2f_WDATA[97] ),
	.h2f_WDATA_98(\arm_a9_hps|fpga_interfaces|h2f_WDATA[98] ),
	.h2f_WDATA_99(\arm_a9_hps|fpga_interfaces|h2f_WDATA[99] ),
	.h2f_WDATA_100(\arm_a9_hps|fpga_interfaces|h2f_WDATA[100] ),
	.h2f_WDATA_101(\arm_a9_hps|fpga_interfaces|h2f_WDATA[101] ),
	.h2f_WDATA_102(\arm_a9_hps|fpga_interfaces|h2f_WDATA[102] ),
	.h2f_WDATA_103(\arm_a9_hps|fpga_interfaces|h2f_WDATA[103] ),
	.h2f_WDATA_104(\arm_a9_hps|fpga_interfaces|h2f_WDATA[104] ),
	.h2f_WDATA_105(\arm_a9_hps|fpga_interfaces|h2f_WDATA[105] ),
	.h2f_WDATA_106(\arm_a9_hps|fpga_interfaces|h2f_WDATA[106] ),
	.h2f_WDATA_107(\arm_a9_hps|fpga_interfaces|h2f_WDATA[107] ),
	.h2f_WDATA_108(\arm_a9_hps|fpga_interfaces|h2f_WDATA[108] ),
	.h2f_WDATA_109(\arm_a9_hps|fpga_interfaces|h2f_WDATA[109] ),
	.h2f_WDATA_110(\arm_a9_hps|fpga_interfaces|h2f_WDATA[110] ),
	.h2f_WDATA_111(\arm_a9_hps|fpga_interfaces|h2f_WDATA[111] ),
	.h2f_WDATA_112(\arm_a9_hps|fpga_interfaces|h2f_WDATA[112] ),
	.h2f_WDATA_113(\arm_a9_hps|fpga_interfaces|h2f_WDATA[113] ),
	.h2f_WDATA_114(\arm_a9_hps|fpga_interfaces|h2f_WDATA[114] ),
	.h2f_WDATA_115(\arm_a9_hps|fpga_interfaces|h2f_WDATA[115] ),
	.h2f_WDATA_116(\arm_a9_hps|fpga_interfaces|h2f_WDATA[116] ),
	.h2f_WDATA_117(\arm_a9_hps|fpga_interfaces|h2f_WDATA[117] ),
	.h2f_WDATA_118(\arm_a9_hps|fpga_interfaces|h2f_WDATA[118] ),
	.h2f_WDATA_119(\arm_a9_hps|fpga_interfaces|h2f_WDATA[119] ),
	.h2f_WDATA_120(\arm_a9_hps|fpga_interfaces|h2f_WDATA[120] ),
	.h2f_WDATA_121(\arm_a9_hps|fpga_interfaces|h2f_WDATA[121] ),
	.h2f_WDATA_122(\arm_a9_hps|fpga_interfaces|h2f_WDATA[122] ),
	.h2f_WDATA_123(\arm_a9_hps|fpga_interfaces|h2f_WDATA[123] ),
	.h2f_WDATA_124(\arm_a9_hps|fpga_interfaces|h2f_WDATA[124] ),
	.h2f_WDATA_125(\arm_a9_hps|fpga_interfaces|h2f_WDATA[125] ),
	.h2f_WDATA_126(\arm_a9_hps|fpga_interfaces|h2f_WDATA[126] ),
	.h2f_WDATA_127(\arm_a9_hps|fpga_interfaces|h2f_WDATA[127] ),
	.h2f_WSTRB_0(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[0] ),
	.h2f_WSTRB_1(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[1] ),
	.h2f_WSTRB_2(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[2] ),
	.h2f_WSTRB_3(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[3] ),
	.h2f_WSTRB_4(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[4] ),
	.h2f_WSTRB_5(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[5] ),
	.h2f_WSTRB_6(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[6] ),
	.h2f_WSTRB_7(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[7] ),
	.h2f_WSTRB_8(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[8] ),
	.h2f_WSTRB_9(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[9] ),
	.h2f_WSTRB_10(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[10] ),
	.h2f_WSTRB_11(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[11] ),
	.h2f_WSTRB_12(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[12] ),
	.h2f_WSTRB_13(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[13] ),
	.h2f_WSTRB_14(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[14] ),
	.h2f_WSTRB_15(\arm_a9_hps|fpga_interfaces|h2f_WSTRB[15] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.sink1_ready(\mm_interconnect_1|cmd_mux|sink1_ready~combout ),
	.awready(\mm_interconnect_1|arm_a9_hps_h2f_lw_axi_master_agent|awready~0_combout ),
	.src0_valid(\mm_interconnect_1|rsp_demux|src0_valid~combout ),
	.source_endofpacket(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent|uncompressor|source_endofpacket~combout ),
	.src1_valid(\mm_interconnect_1|rsp_demux|src1_valid~0_combout ),
	.wready(\mm_interconnect_1|arm_a9_hps_h2f_lw_axi_master_agent|wready~0_combout ),
	.mem_88_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][88]~q ),
	.mem_89_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][89]~q ),
	.mem_90_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][90]~q ),
	.mem_91_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][91]~q ),
	.mem_92_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][99]~q ),
	.out_data_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[0]~0_combout ),
	.out_data_1(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[1]~1_combout ),
	.out_data_2(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[2]~2_combout ),
	.out_data_3(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[3]~3_combout ),
	.out_data_4(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[4]~4_combout ),
	.out_data_5(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[5]~5_combout ),
	.out_data_6(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[6]~6_combout ),
	.out_data_7(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[7]~7_combout ),
	.sink1_ready1(\mm_interconnect_0|cmd_mux_001|sink1_ready~combout ),
	.awready1(\mm_interconnect_0|arm_a9_hps_h2f_axi_master_agent|awready~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.src_payload_0(\mm_interconnect_0|rsp_mux_001|src_payload[0]~combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.wready1(\mm_interconnect_0|arm_a9_hps_h2f_axi_master_agent|wready~0_combout ),
	.src_data_209(\mm_interconnect_0|rsp_mux|src_data[209]~combout ),
	.src_data_210(\mm_interconnect_0|rsp_mux|src_data[210]~combout ),
	.src_data_211(\mm_interconnect_0|rsp_mux|src_data[211]~combout ),
	.src_data_212(\mm_interconnect_0|rsp_mux|src_data[212]~combout ),
	.src_data_213(\mm_interconnect_0|rsp_mux|src_data[213]~combout ),
	.src_data_214(\mm_interconnect_0|rsp_mux|src_data[214]~combout ),
	.src_data_215(\mm_interconnect_0|rsp_mux|src_data[215]~combout ),
	.src_data_216(\mm_interconnect_0|rsp_mux|src_data[216]~combout ),
	.src_data_217(\mm_interconnect_0|rsp_mux|src_data[217]~combout ),
	.src_data_218(\mm_interconnect_0|rsp_mux|src_data[218]~combout ),
	.src_data_219(\mm_interconnect_0|rsp_mux|src_data[219]~combout ),
	.src_data_220(\mm_interconnect_0|rsp_mux|src_data[220]~combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux_001|src_data[0]~1_combout ),
	.src_payload(\mm_interconnect_0|rsp_mux_001|src_payload~4_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux_001|src_data[2]~3_combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux_001|src_data[3]~5_combout ),
	.src_payload1(\mm_interconnect_0|rsp_mux_001|src_payload~6_combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux_001|src_data[5]~7_combout ),
	.src_payload2(\mm_interconnect_0|rsp_mux_001|src_payload~8_combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux_001|src_data[7]~9_combout ),
	.src_payload3(\mm_interconnect_0|rsp_mux_001|src_payload~10_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux_001|src_data[9]~11_combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux_001|src_data[10]~13_combout ),
	.src_data_11(\mm_interconnect_0|rsp_mux_001|src_data[11]~15_combout ),
	.src_data_12(\mm_interconnect_0|rsp_mux_001|src_data[12]~17_combout ),
	.src_payload4(\mm_interconnect_0|rsp_mux_001|src_payload~12_combout ),
	.src_data_14(\mm_interconnect_0|rsp_mux_001|src_data[14]~19_combout ),
	.src_data_15(\mm_interconnect_0|rsp_mux_001|src_data[15]~21_combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux_001|src_data[16]~23_combout ),
	.src_payload5(\mm_interconnect_0|rsp_mux_001|src_payload~14_combout ),
	.src_data_18(\mm_interconnect_0|rsp_mux_001|src_data[18]~25_combout ),
	.src_data_19(\mm_interconnect_0|rsp_mux_001|src_data[19]~27_combout ),
	.src_payload6(\mm_interconnect_0|rsp_mux_001|src_payload~16_combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux_001|src_data[21]~29_combout ),
	.src_payload7(\mm_interconnect_0|rsp_mux_001|src_payload~18_combout ),
	.src_data_23(\mm_interconnect_0|rsp_mux_001|src_data[23]~31_combout ),
	.src_payload8(\mm_interconnect_0|rsp_mux_001|src_payload~20_combout ),
	.src_data_25(\mm_interconnect_0|rsp_mux_001|src_data[25]~33_combout ),
	.src_data_26(\mm_interconnect_0|rsp_mux_001|src_data[26]~35_combout ),
	.src_data_27(\mm_interconnect_0|rsp_mux_001|src_data[27]~37_combout ),
	.src_data_28(\mm_interconnect_0|rsp_mux_001|src_data[28]~39_combout ),
	.src_payload9(\mm_interconnect_0|rsp_mux_001|src_payload~22_combout ),
	.src_data_30(\mm_interconnect_0|rsp_mux_001|src_data[30]~41_combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux_001|src_data[31]~43_combout ),
	.src_data_32(\mm_interconnect_0|rsp_mux_001|src_data[32]~45_combout ),
	.src_payload10(\mm_interconnect_0|rsp_mux_001|src_payload~26_combout ),
	.src_data_34(\mm_interconnect_0|rsp_mux_001|src_data[34]~47_combout ),
	.src_data_35(\mm_interconnect_0|rsp_mux_001|src_data[35]~49_combout ),
	.src_payload11(\mm_interconnect_0|rsp_mux_001|src_payload~28_combout ),
	.src_data_37(\mm_interconnect_0|rsp_mux_001|src_data[37]~51_combout ),
	.src_payload12(\mm_interconnect_0|rsp_mux_001|src_payload~30_combout ),
	.src_data_39(\mm_interconnect_0|rsp_mux_001|src_data[39]~53_combout ),
	.src_payload13(\mm_interconnect_0|rsp_mux_001|src_payload~32_combout ),
	.src_data_41(\mm_interconnect_0|rsp_mux_001|src_data[41]~55_combout ),
	.src_data_42(\mm_interconnect_0|rsp_mux_001|src_data[42]~57_combout ),
	.src_data_43(\mm_interconnect_0|rsp_mux_001|src_data[43]~59_combout ),
	.src_data_44(\mm_interconnect_0|rsp_mux_001|src_data[44]~61_combout ),
	.src_payload14(\mm_interconnect_0|rsp_mux_001|src_payload~34_combout ),
	.src_data_46(\mm_interconnect_0|rsp_mux_001|src_data[46]~63_combout ),
	.src_data_47(\mm_interconnect_0|rsp_mux_001|src_data[47]~65_combout ),
	.src_data_48(\mm_interconnect_0|rsp_mux_001|src_data[48]~67_combout ),
	.src_payload15(\mm_interconnect_0|rsp_mux_001|src_payload~36_combout ),
	.src_data_50(\mm_interconnect_0|rsp_mux_001|src_data[50]~69_combout ),
	.src_data_51(\mm_interconnect_0|rsp_mux_001|src_data[51]~71_combout ),
	.src_payload16(\mm_interconnect_0|rsp_mux_001|src_payload~38_combout ),
	.src_data_53(\mm_interconnect_0|rsp_mux_001|src_data[53]~73_combout ),
	.src_payload17(\mm_interconnect_0|rsp_mux_001|src_payload~40_combout ),
	.src_data_55(\mm_interconnect_0|rsp_mux_001|src_data[55]~75_combout ),
	.src_payload18(\mm_interconnect_0|rsp_mux_001|src_payload~42_combout ),
	.src_data_57(\mm_interconnect_0|rsp_mux_001|src_data[57]~77_combout ),
	.src_data_58(\mm_interconnect_0|rsp_mux_001|src_data[58]~79_combout ),
	.src_data_59(\mm_interconnect_0|rsp_mux_001|src_data[59]~81_combout ),
	.src_data_60(\mm_interconnect_0|rsp_mux_001|src_data[60]~83_combout ),
	.src_payload19(\mm_interconnect_0|rsp_mux_001|src_payload~44_combout ),
	.src_data_62(\mm_interconnect_0|rsp_mux_001|src_data[62]~85_combout ),
	.src_data_63(\mm_interconnect_0|rsp_mux_001|src_data[63]~87_combout ),
	.src_data_64(\mm_interconnect_0|rsp_mux_001|src_data[64]~89_combout ),
	.src_payload20(\mm_interconnect_0|rsp_mux_001|src_payload~48_combout ),
	.src_data_66(\mm_interconnect_0|rsp_mux_001|src_data[66]~91_combout ),
	.src_data_67(\mm_interconnect_0|rsp_mux_001|src_data[67]~93_combout ),
	.src_payload21(\mm_interconnect_0|rsp_mux_001|src_payload~50_combout ),
	.src_data_69(\mm_interconnect_0|rsp_mux_001|src_data[69]~95_combout ),
	.src_payload22(\mm_interconnect_0|rsp_mux_001|src_payload~52_combout ),
	.src_data_71(\mm_interconnect_0|rsp_mux_001|src_data[71]~97_combout ),
	.src_payload23(\mm_interconnect_0|rsp_mux_001|src_payload~54_combout ),
	.src_data_73(\mm_interconnect_0|rsp_mux_001|src_data[73]~99_combout ),
	.src_data_74(\mm_interconnect_0|rsp_mux_001|src_data[74]~101_combout ),
	.src_data_75(\mm_interconnect_0|rsp_mux_001|src_data[75]~103_combout ),
	.src_data_76(\mm_interconnect_0|rsp_mux_001|src_data[76]~105_combout ),
	.src_payload24(\mm_interconnect_0|rsp_mux_001|src_payload~56_combout ),
	.src_data_78(\mm_interconnect_0|rsp_mux_001|src_data[78]~107_combout ),
	.src_data_79(\mm_interconnect_0|rsp_mux_001|src_data[79]~109_combout ),
	.src_data_80(\mm_interconnect_0|rsp_mux_001|src_data[80]~111_combout ),
	.src_payload25(\mm_interconnect_0|rsp_mux_001|src_payload~58_combout ),
	.src_data_82(\mm_interconnect_0|rsp_mux_001|src_data[82]~113_combout ),
	.src_data_83(\mm_interconnect_0|rsp_mux_001|src_data[83]~115_combout ),
	.src_payload26(\mm_interconnect_0|rsp_mux_001|src_payload~60_combout ),
	.src_data_85(\mm_interconnect_0|rsp_mux_001|src_data[85]~117_combout ),
	.src_payload27(\mm_interconnect_0|rsp_mux_001|src_payload~62_combout ),
	.src_data_87(\mm_interconnect_0|rsp_mux_001|src_data[87]~119_combout ),
	.src_payload28(\mm_interconnect_0|rsp_mux_001|src_payload~64_combout ),
	.src_data_89(\mm_interconnect_0|rsp_mux_001|src_data[89]~121_combout ),
	.src_data_90(\mm_interconnect_0|rsp_mux_001|src_data[90]~123_combout ),
	.src_data_91(\mm_interconnect_0|rsp_mux_001|src_data[91]~125_combout ),
	.src_data_92(\mm_interconnect_0|rsp_mux_001|src_data[92]~127_combout ),
	.src_payload29(\mm_interconnect_0|rsp_mux_001|src_payload~66_combout ),
	.src_data_94(\mm_interconnect_0|rsp_mux_001|src_data[94]~129_combout ),
	.src_data_95(\mm_interconnect_0|rsp_mux_001|src_data[95]~131_combout ),
	.src_data_96(\mm_interconnect_0|rsp_mux_001|src_data[96]~combout ),
	.src_payload30(\mm_interconnect_0|rsp_mux_001|src_payload~71_combout ),
	.src_data_98(\mm_interconnect_0|rsp_mux_001|src_data[98]~combout ),
	.src_data_99(\mm_interconnect_0|rsp_mux_001|src_data[99]~combout ),
	.src_payload31(\mm_interconnect_0|rsp_mux_001|src_payload~72_combout ),
	.src_data_101(\mm_interconnect_0|rsp_mux_001|src_data[101]~combout ),
	.src_payload32(\mm_interconnect_0|rsp_mux_001|src_payload~73_combout ),
	.src_data_103(\mm_interconnect_0|rsp_mux_001|src_data[103]~combout ),
	.src_payload33(\mm_interconnect_0|rsp_mux_001|src_payload~74_combout ),
	.src_data_105(\mm_interconnect_0|rsp_mux_001|src_data[105]~combout ),
	.src_data_106(\mm_interconnect_0|rsp_mux_001|src_data[106]~combout ),
	.src_data_107(\mm_interconnect_0|rsp_mux_001|src_data[107]~combout ),
	.src_data_108(\mm_interconnect_0|rsp_mux_001|src_data[108]~combout ),
	.src_payload34(\mm_interconnect_0|rsp_mux_001|src_payload~75_combout ),
	.src_data_110(\mm_interconnect_0|rsp_mux_001|src_data[110]~combout ),
	.src_data_111(\mm_interconnect_0|rsp_mux_001|src_data[111]~combout ),
	.src_data_112(\mm_interconnect_0|rsp_mux_001|src_data[112]~combout ),
	.src_payload35(\mm_interconnect_0|rsp_mux_001|src_payload~76_combout ),
	.src_data_114(\mm_interconnect_0|rsp_mux_001|src_data[114]~combout ),
	.src_data_115(\mm_interconnect_0|rsp_mux_001|src_data[115]~combout ),
	.src_payload36(\mm_interconnect_0|rsp_mux_001|src_payload~77_combout ),
	.src_data_117(\mm_interconnect_0|rsp_mux_001|src_data[117]~combout ),
	.src_payload37(\mm_interconnect_0|rsp_mux_001|src_payload~78_combout ),
	.src_data_119(\mm_interconnect_0|rsp_mux_001|src_data[119]~combout ),
	.src_payload38(\mm_interconnect_0|rsp_mux_001|src_payload~79_combout ),
	.src_data_121(\mm_interconnect_0|rsp_mux_001|src_data[121]~combout ),
	.src_data_122(\mm_interconnect_0|rsp_mux_001|src_data[122]~combout ),
	.src_data_123(\mm_interconnect_0|rsp_mux_001|src_data[123]~combout ),
	.src_data_124(\mm_interconnect_0|rsp_mux_001|src_data[124]~combout ),
	.src_payload39(\mm_interconnect_0|rsp_mux_001|src_payload~80_combout ),
	.src_data_126(\mm_interconnect_0|rsp_mux_001|src_data[126]~combout ),
	.src_data_127(\mm_interconnect_0|rsp_mux_001|src_data[127]~combout ),
	.src_data_2091(\mm_interconnect_0|rsp_mux_001|src_data[209]~combout ),
	.src_data_2101(\mm_interconnect_0|rsp_mux_001|src_data[210]~combout ),
	.src_data_2111(\mm_interconnect_0|rsp_mux_001|src_data[211]~combout ),
	.src_data_2121(\mm_interconnect_0|rsp_mux_001|src_data[212]~combout ),
	.src_data_2131(\mm_interconnect_0|rsp_mux_001|src_data[213]~combout ),
	.src_data_2141(\mm_interconnect_0|rsp_mux_001|src_data[214]~combout ),
	.src_data_2151(\mm_interconnect_0|rsp_mux_001|src_data[215]~combout ),
	.src_data_2161(\mm_interconnect_0|rsp_mux_001|src_data[216]~combout ),
	.src_data_2171(\mm_interconnect_0|rsp_mux_001|src_data[217]~combout ),
	.src_data_2181(\mm_interconnect_0|rsp_mux_001|src_data[218]~combout ),
	.src_data_2191(\mm_interconnect_0|rsp_mux_001|src_data[219]~combout ),
	.src_data_2201(\mm_interconnect_0|rsp_mux_001|src_data[220]~combout ),
	.emac1_inst(\arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_CLK_TX ),
	.emac1_inst1(\arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ),
	.intermediate_0(\arm_a9_hps|hps_io|border|intermediate[0] ),
	.intermediate_1(\arm_a9_hps|hps_io|border|intermediate[1] ),
	.emac1_inst2(\arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ),
	.emac1_inst3(\arm_a9_hps|hps_io|border|emac1_inst~emac_phy_txd ),
	.emac1_inst4(\arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ),
	.emac1_inst5(\arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ),
	.emac1_inst6(\arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ),
	.qspi_inst(\arm_a9_hps|hps_io|border|qspi_inst~O_QSPI_SCLK ),
	.intermediate_2(\arm_a9_hps|hps_io|border|intermediate[2] ),
	.intermediate_4(\arm_a9_hps|hps_io|border|intermediate[4] ),
	.intermediate_6(\arm_a9_hps|hps_io|border|intermediate[6] ),
	.intermediate_8(\arm_a9_hps|hps_io|border|intermediate[8] ),
	.intermediate_3(\arm_a9_hps|hps_io|border|intermediate[3] ),
	.intermediate_5(\arm_a9_hps|hps_io|border|intermediate[5] ),
	.intermediate_7(\arm_a9_hps|hps_io|border|intermediate[7] ),
	.intermediate_9(\arm_a9_hps|hps_io|border|intermediate[9] ),
	.qspi_inst1(\arm_a9_hps|hps_io|border|qspi_inst~O_QSPI_SS_N0 ),
	.sdio_inst(\arm_a9_hps|hps_io|border|sdio_inst~sdmmc_cclk ),
	.intermediate_10(\arm_a9_hps|hps_io|border|intermediate[10] ),
	.intermediate_11(\arm_a9_hps|hps_io|border|intermediate[11] ),
	.intermediate_12(\arm_a9_hps|hps_io|border|intermediate[12] ),
	.intermediate_14(\arm_a9_hps|hps_io|border|intermediate[14] ),
	.intermediate_16(\arm_a9_hps|hps_io|border|intermediate[16] ),
	.intermediate_18(\arm_a9_hps|hps_io|border|intermediate[18] ),
	.intermediate_13(\arm_a9_hps|hps_io|border|intermediate[13] ),
	.intermediate_15(\arm_a9_hps|hps_io|border|intermediate[15] ),
	.intermediate_17(\arm_a9_hps|hps_io|border|intermediate[17] ),
	.intermediate_19(\arm_a9_hps|hps_io|border|intermediate[19] ),
	.usb1_inst(\arm_a9_hps|hps_io|border|usb1_inst~usb_ulpi_stp ),
	.intermediate_20(\arm_a9_hps|hps_io|border|intermediate[20] ),
	.intermediate_22(\arm_a9_hps|hps_io|border|intermediate[22] ),
	.intermediate_24(\arm_a9_hps|hps_io|border|intermediate[24] ),
	.intermediate_26(\arm_a9_hps|hps_io|border|intermediate[26] ),
	.intermediate_28(\arm_a9_hps|hps_io|border|intermediate[28] ),
	.intermediate_30(\arm_a9_hps|hps_io|border|intermediate[30] ),
	.intermediate_32(\arm_a9_hps|hps_io|border|intermediate[32] ),
	.intermediate_34(\arm_a9_hps|hps_io|border|intermediate[34] ),
	.intermediate_21(\arm_a9_hps|hps_io|border|intermediate[21] ),
	.intermediate_23(\arm_a9_hps|hps_io|border|intermediate[23] ),
	.intermediate_25(\arm_a9_hps|hps_io|border|intermediate[25] ),
	.intermediate_27(\arm_a9_hps|hps_io|border|intermediate[27] ),
	.intermediate_29(\arm_a9_hps|hps_io|border|intermediate[29] ),
	.intermediate_31(\arm_a9_hps|hps_io|border|intermediate[31] ),
	.intermediate_33(\arm_a9_hps|hps_io|border|intermediate[33] ),
	.intermediate_35(\arm_a9_hps|hps_io|border|intermediate[35] ),
	.spim1_inst(\arm_a9_hps|hps_io|border|spim1_inst~O_SPI_MASTER_SCLK ),
	.spim1_inst1(\arm_a9_hps|hps_io|border|spim1_inst~O_SPI_MASTER_SS_0_N ),
	.intermediate_36(\arm_a9_hps|hps_io|border|intermediate[36] ),
	.intermediate_37(\arm_a9_hps|hps_io|border|intermediate[37] ),
	.uart0_inst(\arm_a9_hps|hps_io|border|uart0_inst~uart_txd ),
	.intermediate_39(\arm_a9_hps|hps_io|border|intermediate[39] ),
	.intermediate_38(\arm_a9_hps|hps_io|border|intermediate[38] ),
	.intermediate_41(\arm_a9_hps|hps_io|border|intermediate[41] ),
	.intermediate_40(\arm_a9_hps|hps_io|border|intermediate[40] ),
	.intermediate_42(\arm_a9_hps|hps_io|border|intermediate[42] ),
	.intermediate_43(\arm_a9_hps|hps_io|border|intermediate[43] ),
	.intermediate_44(\arm_a9_hps|hps_io|border|intermediate[44] ),
	.intermediate_46(\arm_a9_hps|hps_io|border|intermediate[46] ),
	.intermediate_48(\arm_a9_hps|hps_io|border|intermediate[48] ),
	.intermediate_50(\arm_a9_hps|hps_io|border|intermediate[50] ),
	.intermediate_52(\arm_a9_hps|hps_io|border|intermediate[52] ),
	.intermediate_54(\arm_a9_hps|hps_io|border|intermediate[54] ),
	.intermediate_45(\arm_a9_hps|hps_io|border|intermediate[45] ),
	.intermediate_47(\arm_a9_hps|hps_io|border|intermediate[47] ),
	.intermediate_49(\arm_a9_hps|hps_io|border|intermediate[49] ),
	.intermediate_51(\arm_a9_hps|hps_io|border|intermediate[51] ),
	.intermediate_53(\arm_a9_hps|hps_io|border|intermediate[53] ),
	.intermediate_55(\arm_a9_hps|hps_io|border|intermediate[55] ),
	.intermediate_56(\arm_a9_hps|hps_io|border|intermediate[56] ),
	.intermediate_57(\arm_a9_hps|hps_io|border|intermediate[57] ),
	.parallelterminationcontrol_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] ),
	.parallelterminationcontrol_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ),
	.parallelterminationcontrol_2(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ),
	.parallelterminationcontrol_3(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ),
	.parallelterminationcontrol_4(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ),
	.parallelterminationcontrol_5(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ),
	.parallelterminationcontrol_6(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ),
	.parallelterminationcontrol_7(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ),
	.parallelterminationcontrol_8(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ),
	.parallelterminationcontrol_9(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ),
	.parallelterminationcontrol_10(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ),
	.parallelterminationcontrol_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ),
	.parallelterminationcontrol_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ),
	.parallelterminationcontrol_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ),
	.parallelterminationcontrol_14(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ),
	.parallelterminationcontrol_15(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ),
	.seriesterminationcontrol_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] ),
	.seriesterminationcontrol_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ),
	.seriesterminationcontrol_2(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ),
	.seriesterminationcontrol_3(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ),
	.seriesterminationcontrol_4(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ),
	.seriesterminationcontrol_5(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ),
	.seriesterminationcontrol_6(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ),
	.seriesterminationcontrol_7(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ),
	.seriesterminationcontrol_8(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ),
	.seriesterminationcontrol_9(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ),
	.seriesterminationcontrol_10(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ),
	.seriesterminationcontrol_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ),
	.seriesterminationcontrol_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ),
	.seriesterminationcontrol_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ),
	.seriesterminationcontrol_14(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ),
	.seriesterminationcontrol_15(\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ),
	.dqsin(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dataout_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ),
	.dataout_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ),
	.dataout_2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ),
	.dataout_3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ),
	.dataout_4(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ),
	.dataout_5(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ),
	.dataout_6(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ),
	.dataout_7(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ),
	.dataout_8(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ),
	.dataout_9(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ),
	.dataout_10(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ),
	.dataout_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ),
	.dataout_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ),
	.dataout_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ),
	.dataout_14(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ),
	.dataout_01(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ),
	.dataout_15(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ),
	.dataout_21(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ),
	.dataout_16(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ),
	.dataout_02(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ),
	.dataout_31(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ),
	.dataout_41(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ),
	.dataout_51(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ),
	.dataout_03(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ),
	.dataout_22(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ),
	.extra_output_pad_gen0delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.wire_pseudo_diffa_o_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ),
	.wire_pseudo_diffa_obar_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ),
	.wire_pseudo_diffa_oeout_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ),
	.wire_pseudo_diffa_oebout_0(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ),
	.pad_gen0delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_11(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_12(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_13(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.os(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar1(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar2(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar3(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.hps_io_emac1_inst_MDIO_0(\arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o ),
	.hps_io_qspi_inst_IO0_0(\arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~input_o ),
	.hps_io_qspi_inst_IO1_0(\arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~input_o ),
	.hps_io_qspi_inst_IO2_0(\arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~input_o ),
	.hps_io_qspi_inst_IO3_0(\arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~input_o ),
	.hps_io_sdio_inst_CMD_0(\arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o ),
	.hps_io_sdio_inst_D0_0(\arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~input_o ),
	.hps_io_sdio_inst_D1_0(\arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~input_o ),
	.hps_io_sdio_inst_D2_0(\arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~input_o ),
	.hps_io_sdio_inst_D3_0(\arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~input_o ),
	.hps_io_usb1_inst_D0_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~input_o ),
	.hps_io_usb1_inst_D1_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~input_o ),
	.hps_io_usb1_inst_D2_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~input_o ),
	.hps_io_usb1_inst_D3_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~input_o ),
	.hps_io_usb1_inst_D4_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~input_o ),
	.hps_io_usb1_inst_D5_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~input_o ),
	.hps_io_usb1_inst_D6_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~input_o ),
	.hps_io_usb1_inst_D7_0(\arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~input_o ),
	.hps_io_i2c0_inst_SDA_0(\arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~input_o ),
	.hps_io_i2c0_inst_SCL_0(\arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~input_o ),
	.hps_io_i2c1_inst_SDA_0(\arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~input_o ),
	.hps_io_i2c1_inst_SCL_0(\arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~input_o ),
	.hps_io_gpio_inst_GPIO09_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~input_o ),
	.hps_io_gpio_inst_GPIO35_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~input_o ),
	.hps_io_gpio_inst_GPIO40_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~input_o ),
	.hps_io_gpio_inst_GPIO41_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~input_o ),
	.hps_io_gpio_inst_GPIO48_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~input_o ),
	.hps_io_gpio_inst_GPIO53_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~input_o ),
	.hps_io_gpio_inst_GPIO54_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~input_o ),
	.hps_io_gpio_inst_GPIO61_0(\arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~input_o ),
	.hps_io_hps_io_emac1_inst_RXD0(\hps_io_hps_io_emac1_inst_RXD0~input_o ),
	.hps_io_hps_io_emac1_inst_RXD1(\hps_io_hps_io_emac1_inst_RXD1~input_o ),
	.hps_io_hps_io_emac1_inst_RXD2(\hps_io_hps_io_emac1_inst_RXD2~input_o ),
	.hps_io_hps_io_emac1_inst_RXD3(\hps_io_hps_io_emac1_inst_RXD3~input_o ),
	.hps_io_hps_io_emac1_inst_RX_CLK(\hps_io_hps_io_emac1_inst_RX_CLK~input_o ),
	.hps_io_hps_io_emac1_inst_RX_CTL(\hps_io_hps_io_emac1_inst_RX_CTL~input_o ),
	.hps_io_hps_io_spim1_inst_MISO(\hps_io_hps_io_spim1_inst_MISO~input_o ),
	.hps_io_hps_io_uart0_inst_RX(\hps_io_hps_io_uart0_inst_RX~input_o ),
	.hps_io_hps_io_usb1_inst_CLK(\hps_io_hps_io_usb1_inst_CLK~input_o ),
	.hps_io_hps_io_usb1_inst_DIR(\hps_io_hps_io_usb1_inst_DIR~input_o ),
	.hps_io_hps_io_usb1_inst_NXT(\hps_io_hps_io_usb1_inst_NXT~input_o ),
	.memory_oct_rzqin(\memory_oct_rzqin~input_o ));

Computer_System_altera_reset_controller_2 rst_controller_002(
	.h2f_rst_n_0(\arm_a9_hps|fpga_interfaces|h2f_rst_n[0] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ));

Computer_System_altera_reset_controller_1 rst_controller_001(
	.h2f_rst_n_0(\arm_a9_hps|fpga_interfaces|h2f_rst_n[0] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.locked_wire_0(\system_pll|sys_pll|altera_pll_i|locked_wire[0] ),
	.r_early_rst1(\rst_controller_001|r_early_rst~q ),
	.r_sync_rst1(\rst_controller_001|r_sync_rst~q ),
	.merged_reset(\rst_controller_001|merged_reset~0_combout ));

Computer_System_altera_reset_controller rst_controller(
	.r_sync_rst1(\rst_controller|r_sync_rst~q ),
	.r_early_rst1(\rst_controller|r_early_rst~q ),
	.merged_reset(\rst_controller_001|merged_reset~0_combout ),
	.clock_bridge_0_in_clk_clk(\clock_bridge_0_in_clk_clk~input_o ));

Computer_System_Computer_System_mm_interconnect_1 mm_interconnect_1(
	.h2f_lw_ARVALID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARVALID[0] ),
	.h2f_lw_AWVALID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWVALID[0] ),
	.h2f_lw_BREADY_0(\arm_a9_hps|fpga_interfaces|h2f_lw_BREADY[0] ),
	.h2f_lw_RREADY_0(\arm_a9_hps|fpga_interfaces|h2f_lw_RREADY[0] ),
	.h2f_lw_WLAST_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WLAST[0] ),
	.h2f_lw_WVALID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WVALID[0] ),
	.h2f_lw_ARADDR_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[0] ),
	.h2f_lw_ARADDR_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[1] ),
	.h2f_lw_ARADDR_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[2] ),
	.h2f_lw_ARADDR_3(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[3] ),
	.h2f_lw_ARADDR_4(\arm_a9_hps|fpga_interfaces|h2f_lw_ARADDR[4] ),
	.h2f_lw_ARBURST_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARBURST[0] ),
	.h2f_lw_ARBURST_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARBURST[1] ),
	.h2f_lw_ARID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[0] ),
	.h2f_lw_ARID_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[1] ),
	.h2f_lw_ARID_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[2] ),
	.h2f_lw_ARID_3(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[3] ),
	.h2f_lw_ARID_4(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[4] ),
	.h2f_lw_ARID_5(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[5] ),
	.h2f_lw_ARID_6(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[6] ),
	.h2f_lw_ARID_7(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[7] ),
	.h2f_lw_ARID_8(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[8] ),
	.h2f_lw_ARID_9(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[9] ),
	.h2f_lw_ARID_10(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[10] ),
	.h2f_lw_ARID_11(\arm_a9_hps|fpga_interfaces|h2f_lw_ARID[11] ),
	.h2f_lw_ARLEN_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[0] ),
	.h2f_lw_ARLEN_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[1] ),
	.h2f_lw_ARLEN_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[2] ),
	.h2f_lw_ARLEN_3(\arm_a9_hps|fpga_interfaces|h2f_lw_ARLEN[3] ),
	.h2f_lw_ARSIZE_0(\arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[0] ),
	.h2f_lw_ARSIZE_1(\arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[1] ),
	.h2f_lw_ARSIZE_2(\arm_a9_hps|fpga_interfaces|h2f_lw_ARSIZE[2] ),
	.h2f_lw_AWADDR_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[0] ),
	.h2f_lw_AWADDR_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[1] ),
	.h2f_lw_AWADDR_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[2] ),
	.h2f_lw_AWADDR_3(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[3] ),
	.h2f_lw_AWADDR_4(\arm_a9_hps|fpga_interfaces|h2f_lw_AWADDR[4] ),
	.h2f_lw_AWBURST_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWBURST[0] ),
	.h2f_lw_AWBURST_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWBURST[1] ),
	.h2f_lw_AWID_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[0] ),
	.h2f_lw_AWID_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[1] ),
	.h2f_lw_AWID_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[2] ),
	.h2f_lw_AWID_3(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[3] ),
	.h2f_lw_AWID_4(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[4] ),
	.h2f_lw_AWID_5(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[5] ),
	.h2f_lw_AWID_6(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[6] ),
	.h2f_lw_AWID_7(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[7] ),
	.h2f_lw_AWID_8(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[8] ),
	.h2f_lw_AWID_9(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[9] ),
	.h2f_lw_AWID_10(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[10] ),
	.h2f_lw_AWID_11(\arm_a9_hps|fpga_interfaces|h2f_lw_AWID[11] ),
	.h2f_lw_AWLEN_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[0] ),
	.h2f_lw_AWLEN_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[1] ),
	.h2f_lw_AWLEN_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[2] ),
	.h2f_lw_AWLEN_3(\arm_a9_hps|fpga_interfaces|h2f_lw_AWLEN[3] ),
	.h2f_lw_AWSIZE_0(\arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[0] ),
	.h2f_lw_AWSIZE_1(\arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[1] ),
	.h2f_lw_AWSIZE_2(\arm_a9_hps|fpga_interfaces|h2f_lw_AWSIZE[2] ),
	.h2f_lw_WDATA_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[0] ),
	.h2f_lw_WDATA_1(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[1] ),
	.h2f_lw_WDATA_2(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[2] ),
	.h2f_lw_WDATA_3(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[3] ),
	.h2f_lw_WDATA_4(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[4] ),
	.h2f_lw_WDATA_5(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[5] ),
	.h2f_lw_WDATA_6(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[6] ),
	.h2f_lw_WDATA_7(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[7] ),
	.h2f_lw_WDATA_8(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[8] ),
	.h2f_lw_WDATA_9(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[9] ),
	.h2f_lw_WDATA_10(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[10] ),
	.h2f_lw_WDATA_11(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[11] ),
	.h2f_lw_WDATA_12(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[12] ),
	.h2f_lw_WDATA_13(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[13] ),
	.h2f_lw_WDATA_14(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[14] ),
	.h2f_lw_WDATA_15(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[15] ),
	.h2f_lw_WDATA_16(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[16] ),
	.h2f_lw_WDATA_17(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[17] ),
	.h2f_lw_WDATA_18(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[18] ),
	.h2f_lw_WDATA_19(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[19] ),
	.h2f_lw_WDATA_20(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[20] ),
	.h2f_lw_WDATA_21(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[21] ),
	.h2f_lw_WDATA_22(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[22] ),
	.h2f_lw_WDATA_23(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[23] ),
	.h2f_lw_WDATA_24(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[24] ),
	.h2f_lw_WDATA_25(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[25] ),
	.h2f_lw_WDATA_26(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[26] ),
	.h2f_lw_WDATA_27(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[27] ),
	.h2f_lw_WDATA_28(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[28] ),
	.h2f_lw_WDATA_29(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[29] ),
	.h2f_lw_WDATA_30(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[30] ),
	.h2f_lw_WDATA_31(\arm_a9_hps|fpga_interfaces|h2f_lw_WDATA[31] ),
	.h2f_lw_WSTRB_0(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[0] ),
	.h2f_lw_WSTRB_1(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[1] ),
	.h2f_lw_WSTRB_2(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[2] ),
	.h2f_lw_WSTRB_3(\arm_a9_hps|fpga_interfaces|h2f_lw_WSTRB[3] ),
	.outclk_wire_0(\system_pll|sys_pll|altera_pll_i|outclk_wire[0] ),
	.in_ready_hold(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.wait_latency_counter_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_1(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_translator|wait_latency_counter[1]~q ),
	.sink1_ready(\mm_interconnect_1|cmd_mux|sink1_ready~combout ),
	.ARM_A9_HPS_h2f_lw_axi_master_awready(\mm_interconnect_1|arm_a9_hps_h2f_lw_axi_master_agent|awready~0_combout ),
	.src0_valid(\mm_interconnect_1|rsp_demux|src0_valid~combout ),
	.source_endofpacket(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent|uncompressor|source_endofpacket~combout ),
	.src1_valid(\mm_interconnect_1|rsp_demux|src1_valid~0_combout ),
	.ARM_A9_HPS_h2f_lw_axi_master_wready(\mm_interconnect_1|arm_a9_hps_h2f_lw_axi_master_agent|wready~0_combout ),
	.mem_88_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][88]~q ),
	.mem_89_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][89]~q ),
	.mem_90_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][90]~q ),
	.mem_91_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][91]~q ),
	.mem_92_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][99]~q ),
	.out_data_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[0]~0_combout ),
	.out_data_1(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[1]~1_combout ),
	.out_data_2(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[2]~2_combout ),
	.out_data_3(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[3]~3_combout ),
	.out_data_4(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[4]~4_combout ),
	.out_data_5(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[5]~5_combout ),
	.out_data_6(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[6]~6_combout ),
	.out_data_7(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent_rdata_fifo|out_data[7]~7_combout ),
	.r_sync_rst(\rst_controller_001|r_sync_rst~q ),
	.m0_write(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent|m0_write~combout ),
	.m0_read(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_agent|m0_read~0_combout ),
	.wrclk_control_slave_readdata_0(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[0]~q ),
	.wrclk_control_slave_readdata_1(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[1]~q ),
	.wrclk_control_slave_readdata_2(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[2]~q ),
	.wrclk_control_slave_readdata_3(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[3]~q ),
	.wrclk_control_slave_readdata_4(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[4]~q ),
	.wrclk_control_slave_readdata_5(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[5]~q ),
	.wrclk_control_slave_readdata_6(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[6]~q ),
	.wrclk_control_slave_readdata_7(\fifo_hps_to_fpga|the_dcfifo_with_controls|wrclk_control_slave_readdata[7]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_002|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_4(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[4]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.in_data_reg_0(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.in_data_reg_2(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_1(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_14(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_8(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_13(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_12(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_11(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_10(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_9(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_19(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_18(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_17(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_16(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_15(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_26(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_21(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_20(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_31(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.in_data_reg_30(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_29(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_28(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_27(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_25(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_24(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.in_data_reg_23(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_22(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_7(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_6(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_5(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_4(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_3(\mm_interconnect_1|fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ));

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[3]),
	.ibar(memory_mem_dqs_n[3]),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[24]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[25]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[26]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[27]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[28]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[29]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[30]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[31]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[2]),
	.ibar(memory_mem_dqs_n[2]),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[16]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[17]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[18]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[19]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[20]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[21]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[22]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[23]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[1]),
	.ibar(memory_mem_dqs_n[1]),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[8]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[9]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[10]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[11]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[12]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[13]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[14]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[15]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[0]),
	.ibar(memory_mem_dqs_n[0]),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[0]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[1]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[2]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[3]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[4]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[5]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[6]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[7]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

assign \arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o  = hps_io_hps_io_emac1_inst_MDIO;

assign \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~input_o  = hps_io_hps_io_qspi_inst_IO0;

assign \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~input_o  = hps_io_hps_io_qspi_inst_IO1;

assign \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~input_o  = hps_io_hps_io_qspi_inst_IO2;

assign \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~input_o  = hps_io_hps_io_qspi_inst_IO3;

assign \arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o  = hps_io_hps_io_sdio_inst_CMD;

assign \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~input_o  = hps_io_hps_io_sdio_inst_D0;

assign \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~input_o  = hps_io_hps_io_sdio_inst_D1;

assign \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~input_o  = hps_io_hps_io_sdio_inst_D2;

assign \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~input_o  = hps_io_hps_io_sdio_inst_D3;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~input_o  = hps_io_hps_io_usb1_inst_D0;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~input_o  = hps_io_hps_io_usb1_inst_D1;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~input_o  = hps_io_hps_io_usb1_inst_D2;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~input_o  = hps_io_hps_io_usb1_inst_D3;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~input_o  = hps_io_hps_io_usb1_inst_D4;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~input_o  = hps_io_hps_io_usb1_inst_D5;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~input_o  = hps_io_hps_io_usb1_inst_D6;

assign \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~input_o  = hps_io_hps_io_usb1_inst_D7;

assign \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~input_o  = hps_io_hps_io_i2c0_inst_SDA;

assign \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~input_o  = hps_io_hps_io_i2c0_inst_SCL;

assign \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~input_o  = hps_io_hps_io_i2c1_inst_SDA;

assign \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~input_o  = hps_io_hps_io_i2c1_inst_SCL;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO09;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO35;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO40;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO41;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO48;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO53;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO54;

assign \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~input_o  = hps_io_hps_io_gpio_inst_GPIO61;

assign \hps_io_hps_io_emac1_inst_RXD0~input_o  = hps_io_hps_io_emac1_inst_RXD0;

assign \hps_io_hps_io_emac1_inst_RXD1~input_o  = hps_io_hps_io_emac1_inst_RXD1;

assign \hps_io_hps_io_emac1_inst_RXD2~input_o  = hps_io_hps_io_emac1_inst_RXD2;

assign \hps_io_hps_io_emac1_inst_RXD3~input_o  = hps_io_hps_io_emac1_inst_RXD3;

assign \hps_io_hps_io_emac1_inst_RX_CLK~input_o  = hps_io_hps_io_emac1_inst_RX_CLK;

assign \hps_io_hps_io_emac1_inst_RX_CTL~input_o  = hps_io_hps_io_emac1_inst_RX_CTL;

assign \hps_io_hps_io_spim1_inst_MISO~input_o  = hps_io_hps_io_spim1_inst_MISO;

assign \hps_io_hps_io_uart0_inst_RX~input_o  = hps_io_hps_io_uart0_inst_RX;

assign \hps_io_hps_io_usb1_inst_CLK~input_o  = hps_io_hps_io_usb1_inst_CLK;

assign \hps_io_hps_io_usb1_inst_DIR~input_o  = hps_io_hps_io_usb1_inst_DIR;

assign \hps_io_hps_io_usb1_inst_NXT~input_o  = hps_io_hps_io_usb1_inst_NXT;

assign \memory_oct_rzqin~input_o  = memory_oct_rzqin;

assign \fifo_hps_to_fpga_out_read~input_o  = fifo_hps_to_fpga_out_read;

assign \clock_bridge_0_in_clk_clk~input_o  = clock_bridge_0_in_clk_clk;

assign \fifo_hps_to_fpga_out_csr_address[2]~input_o  = fifo_hps_to_fpga_out_csr_address[2];

assign \fifo_hps_to_fpga_out_csr_address[0]~input_o  = fifo_hps_to_fpga_out_csr_address[0];

assign \fifo_hps_to_fpga_out_csr_address[1]~input_o  = fifo_hps_to_fpga_out_csr_address[1];

assign \fifo_hps_to_fpga_out_csr_read~input_o  = fifo_hps_to_fpga_out_csr_read;

assign \onchip_sram_s1_chipselect~input_o  = onchip_sram_s1_chipselect;

assign \onchip_sram_s1_write~input_o  = onchip_sram_s1_write;

assign \onchip_sram_s1_clken~input_o  = onchip_sram_s1_clken;

assign \onchip_sram_s1_writedata[0]~input_o  = onchip_sram_s1_writedata[0];

assign \onchip_sram_s1_address[0]~input_o  = onchip_sram_s1_address[0];

assign \onchip_sram_s1_address[1]~input_o  = onchip_sram_s1_address[1];

assign \onchip_sram_s1_address[2]~input_o  = onchip_sram_s1_address[2];

assign \onchip_sram_s1_address[3]~input_o  = onchip_sram_s1_address[3];

assign \onchip_sram_s1_address[4]~input_o  = onchip_sram_s1_address[4];

assign \onchip_sram_s1_address[5]~input_o  = onchip_sram_s1_address[5];

assign \onchip_sram_s1_address[6]~input_o  = onchip_sram_s1_address[6];

assign \onchip_sram_s1_address[7]~input_o  = onchip_sram_s1_address[7];

assign \onchip_sram_s1_byteenable[0]~input_o  = onchip_sram_s1_byteenable[0];

assign \onchip_sram_s1_writedata[1]~input_o  = onchip_sram_s1_writedata[1];

assign \onchip_sram_s1_writedata[2]~input_o  = onchip_sram_s1_writedata[2];

assign \onchip_sram_s1_writedata[3]~input_o  = onchip_sram_s1_writedata[3];

assign \onchip_sram_s1_writedata[4]~input_o  = onchip_sram_s1_writedata[4];

assign \onchip_sram_s1_writedata[5]~input_o  = onchip_sram_s1_writedata[5];

assign \onchip_sram_s1_writedata[6]~input_o  = onchip_sram_s1_writedata[6];

assign \onchip_sram_s1_writedata[7]~input_o  = onchip_sram_s1_writedata[7];

assign \onchip_sram_s1_writedata[8]~input_o  = onchip_sram_s1_writedata[8];

assign \onchip_sram_s1_byteenable[1]~input_o  = onchip_sram_s1_byteenable[1];

assign \onchip_sram_s1_writedata[9]~input_o  = onchip_sram_s1_writedata[9];

assign \onchip_sram_s1_writedata[10]~input_o  = onchip_sram_s1_writedata[10];

assign \onchip_sram_s1_writedata[11]~input_o  = onchip_sram_s1_writedata[11];

assign \onchip_sram_s1_writedata[12]~input_o  = onchip_sram_s1_writedata[12];

assign \onchip_sram_s1_writedata[13]~input_o  = onchip_sram_s1_writedata[13];

assign \onchip_sram_s1_writedata[14]~input_o  = onchip_sram_s1_writedata[14];

assign \onchip_sram_s1_writedata[15]~input_o  = onchip_sram_s1_writedata[15];

assign \onchip_sram_s1_writedata[16]~input_o  = onchip_sram_s1_writedata[16];

assign \onchip_sram_s1_byteenable[2]~input_o  = onchip_sram_s1_byteenable[2];

assign \onchip_sram_s1_writedata[17]~input_o  = onchip_sram_s1_writedata[17];

assign \onchip_sram_s1_writedata[18]~input_o  = onchip_sram_s1_writedata[18];

assign \onchip_sram_s1_writedata[19]~input_o  = onchip_sram_s1_writedata[19];

assign \onchip_sram_s1_writedata[20]~input_o  = onchip_sram_s1_writedata[20];

assign \onchip_sram_s1_writedata[21]~input_o  = onchip_sram_s1_writedata[21];

assign \onchip_sram_s1_writedata[22]~input_o  = onchip_sram_s1_writedata[22];

assign \onchip_sram_s1_writedata[23]~input_o  = onchip_sram_s1_writedata[23];

assign \onchip_sram_s1_writedata[24]~input_o  = onchip_sram_s1_writedata[24];

assign \onchip_sram_s1_byteenable[3]~input_o  = onchip_sram_s1_byteenable[3];

assign \onchip_sram_s1_writedata[25]~input_o  = onchip_sram_s1_writedata[25];

assign \onchip_sram_s1_writedata[26]~input_o  = onchip_sram_s1_writedata[26];

assign \onchip_sram_s1_writedata[27]~input_o  = onchip_sram_s1_writedata[27];

assign \onchip_sram_s1_writedata[28]~input_o  = onchip_sram_s1_writedata[28];

assign \onchip_sram_s1_writedata[29]~input_o  = onchip_sram_s1_writedata[29];

assign \onchip_sram_s1_writedata[30]~input_o  = onchip_sram_s1_writedata[30];

assign \onchip_sram_s1_writedata[31]~input_o  = onchip_sram_s1_writedata[31];

assign \system_pll_ref_clk_clk~input_o  = system_pll_ref_clk_clk;

assign \system_pll_ref_reset_reset~input_o  = system_pll_ref_reset_reset;

assign \fifo_hps_to_fpga_out_csr_writedata[0]~input_o  = fifo_hps_to_fpga_out_csr_writedata[0];

assign \fifo_hps_to_fpga_out_csr_write~input_o  = fifo_hps_to_fpga_out_csr_write;

assign \fifo_hps_to_fpga_out_csr_writedata[7]~input_o  = fifo_hps_to_fpga_out_csr_writedata[7];

assign \fifo_hps_to_fpga_out_csr_writedata[1]~input_o  = fifo_hps_to_fpga_out_csr_writedata[1];

assign \fifo_hps_to_fpga_out_csr_writedata[13]~input_o  = fifo_hps_to_fpga_out_csr_writedata[13];

assign \fifo_hps_to_fpga_out_csr_writedata[19]~input_o  = fifo_hps_to_fpga_out_csr_writedata[19];

assign \fifo_hps_to_fpga_out_csr_writedata[26]~input_o  = fifo_hps_to_fpga_out_csr_writedata[26];

assign \fifo_hps_to_fpga_out_csr_writedata[27]~input_o  = fifo_hps_to_fpga_out_csr_writedata[27];

assign \fifo_hps_to_fpga_out_csr_writedata[28]~input_o  = fifo_hps_to_fpga_out_csr_writedata[28];

assign \fifo_hps_to_fpga_out_csr_writedata[29]~input_o  = fifo_hps_to_fpga_out_csr_writedata[29];

assign \fifo_hps_to_fpga_out_csr_writedata[30]~input_o  = fifo_hps_to_fpga_out_csr_writedata[30];

assign \fifo_hps_to_fpga_out_csr_writedata[31]~input_o  = fifo_hps_to_fpga_out_csr_writedata[31];

assign \fifo_hps_to_fpga_out_csr_writedata[20]~input_o  = fifo_hps_to_fpga_out_csr_writedata[20];

assign \fifo_hps_to_fpga_out_csr_writedata[21]~input_o  = fifo_hps_to_fpga_out_csr_writedata[21];

assign \fifo_hps_to_fpga_out_csr_writedata[22]~input_o  = fifo_hps_to_fpga_out_csr_writedata[22];

assign \fifo_hps_to_fpga_out_csr_writedata[23]~input_o  = fifo_hps_to_fpga_out_csr_writedata[23];

assign \fifo_hps_to_fpga_out_csr_writedata[24]~input_o  = fifo_hps_to_fpga_out_csr_writedata[24];

assign \fifo_hps_to_fpga_out_csr_writedata[25]~input_o  = fifo_hps_to_fpga_out_csr_writedata[25];

assign \fifo_hps_to_fpga_out_csr_writedata[8]~input_o  = fifo_hps_to_fpga_out_csr_writedata[8];

assign \fifo_hps_to_fpga_out_csr_writedata[9]~input_o  = fifo_hps_to_fpga_out_csr_writedata[9];

assign \fifo_hps_to_fpga_out_csr_writedata[10]~input_o  = fifo_hps_to_fpga_out_csr_writedata[10];

assign \fifo_hps_to_fpga_out_csr_writedata[11]~input_o  = fifo_hps_to_fpga_out_csr_writedata[11];

assign \fifo_hps_to_fpga_out_csr_writedata[12]~input_o  = fifo_hps_to_fpga_out_csr_writedata[12];

assign \fifo_hps_to_fpga_out_csr_writedata[14]~input_o  = fifo_hps_to_fpga_out_csr_writedata[14];

assign \fifo_hps_to_fpga_out_csr_writedata[15]~input_o  = fifo_hps_to_fpga_out_csr_writedata[15];

assign \fifo_hps_to_fpga_out_csr_writedata[16]~input_o  = fifo_hps_to_fpga_out_csr_writedata[16];

assign \fifo_hps_to_fpga_out_csr_writedata[17]~input_o  = fifo_hps_to_fpga_out_csr_writedata[17];

assign \fifo_hps_to_fpga_out_csr_writedata[18]~input_o  = fifo_hps_to_fpga_out_csr_writedata[18];

assign \fifo_hps_to_fpga_out_csr_writedata[2]~input_o  = fifo_hps_to_fpga_out_csr_writedata[2];

assign \fifo_hps_to_fpga_out_csr_writedata[3]~input_o  = fifo_hps_to_fpga_out_csr_writedata[3];

assign \fifo_hps_to_fpga_out_csr_writedata[4]~input_o  = fifo_hps_to_fpga_out_csr_writedata[4];

assign \fifo_hps_to_fpga_out_csr_writedata[5]~input_o  = fifo_hps_to_fpga_out_csr_writedata[5];

assign \fifo_hps_to_fpga_out_csr_writedata[6]~input_o  = fifo_hps_to_fpga_out_csr_writedata[6];

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[3]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[2]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[1]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[0]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(memory_mem_ck_n),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(memory_mem_ck),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_spim1_inst_MOSI[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[36] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[37] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_spim1_inst_MOSI),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_spim1_inst_MOSI[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_spim1_inst_MOSI[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_spim1_inst_MOSI[0]~output .shift_series_termination_control = "false";

assign fifo_hps_to_fpga_out_readdata[0] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[0] ;

assign fifo_hps_to_fpga_out_readdata[1] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[1] ;

assign fifo_hps_to_fpga_out_readdata[2] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[2] ;

assign fifo_hps_to_fpga_out_readdata[3] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[3] ;

assign fifo_hps_to_fpga_out_readdata[4] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[4] ;

assign fifo_hps_to_fpga_out_readdata[5] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[5] ;

assign fifo_hps_to_fpga_out_readdata[6] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[6] ;

assign fifo_hps_to_fpga_out_readdata[7] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[7] ;

assign fifo_hps_to_fpga_out_readdata[8] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[8] ;

assign fifo_hps_to_fpga_out_readdata[9] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[9] ;

assign fifo_hps_to_fpga_out_readdata[10] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[10] ;

assign fifo_hps_to_fpga_out_readdata[11] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[11] ;

assign fifo_hps_to_fpga_out_readdata[12] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[12] ;

assign fifo_hps_to_fpga_out_readdata[13] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[13] ;

assign fifo_hps_to_fpga_out_readdata[14] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[14] ;

assign fifo_hps_to_fpga_out_readdata[15] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[15] ;

assign fifo_hps_to_fpga_out_readdata[16] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[16] ;

assign fifo_hps_to_fpga_out_readdata[17] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[17] ;

assign fifo_hps_to_fpga_out_readdata[18] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[18] ;

assign fifo_hps_to_fpga_out_readdata[19] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[19] ;

assign fifo_hps_to_fpga_out_readdata[20] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[20] ;

assign fifo_hps_to_fpga_out_readdata[21] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[21] ;

assign fifo_hps_to_fpga_out_readdata[22] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[22] ;

assign fifo_hps_to_fpga_out_readdata[23] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[23] ;

assign fifo_hps_to_fpga_out_readdata[24] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[24] ;

assign fifo_hps_to_fpga_out_readdata[25] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[25] ;

assign fifo_hps_to_fpga_out_readdata[26] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[26] ;

assign fifo_hps_to_fpga_out_readdata[27] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[27] ;

assign fifo_hps_to_fpga_out_readdata[28] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[28] ;

assign fifo_hps_to_fpga_out_readdata[29] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[29] ;

assign fifo_hps_to_fpga_out_readdata[30] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[30] ;

assign fifo_hps_to_fpga_out_readdata[31] = \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|fifo_ram|q_b[31] ;

assign fifo_hps_to_fpga_out_waitrequest = ~ \fifo_hps_to_fpga|the_dcfifo_with_controls|the_dcfifo|dual_clock_fifo|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~combout ;

assign fifo_hps_to_fpga_out_csr_readdata[0] = \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[0]~q ;

assign fifo_hps_to_fpga_out_csr_readdata[1] = \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[1]~q ;

assign fifo_hps_to_fpga_out_csr_readdata[2] = \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[2]~q ;

assign fifo_hps_to_fpga_out_csr_readdata[3] = \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[3]~q ;

assign fifo_hps_to_fpga_out_csr_readdata[4] = \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[4]~q ;

assign fifo_hps_to_fpga_out_csr_readdata[5] = \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[5]~q ;

assign fifo_hps_to_fpga_out_csr_readdata[6] = \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[6]~q ;

assign fifo_hps_to_fpga_out_csr_readdata[7] = \fifo_hps_to_fpga|the_dcfifo_with_controls|rdclk_control_slave_readdata[7]~q ;

assign fifo_hps_to_fpga_out_csr_readdata[8] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[9] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[10] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[11] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[12] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[13] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[14] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[15] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[16] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[17] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[18] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[19] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[20] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[21] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[22] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[23] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[24] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[25] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[26] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[27] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[28] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[29] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[30] = gnd;

assign fifo_hps_to_fpga_out_csr_readdata[31] = gnd;

assign hps_io_hps_io_emac1_inst_TX_CLK = \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_CLK_TX ;

assign hps_io_hps_io_emac1_inst_TXD0 = \arm_a9_hps|hps_io|border|emac1_inst~emac_phy_txd ;

assign hps_io_hps_io_emac1_inst_TXD1 = \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ;

assign hps_io_hps_io_emac1_inst_TXD2 = \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ;

assign hps_io_hps_io_emac1_inst_TXD3 = \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ;

assign hps_io_hps_io_emac1_inst_MDC = \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ;

assign hps_io_hps_io_emac1_inst_TX_CTL = \arm_a9_hps|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ;

assign hps_io_hps_io_qspi_inst_SS0 = \arm_a9_hps|hps_io|border|qspi_inst~O_QSPI_SS_N0 ;

assign hps_io_hps_io_qspi_inst_CLK = \arm_a9_hps|hps_io|border|qspi_inst~O_QSPI_SCLK ;

assign hps_io_hps_io_sdio_inst_CLK = \arm_a9_hps|hps_io|border|sdio_inst~sdmmc_cclk ;

assign hps_io_hps_io_usb1_inst_STP = \arm_a9_hps|hps_io|border|usb1_inst~usb_ulpi_stp ;

assign hps_io_hps_io_spim1_inst_CLK = \arm_a9_hps|hps_io|border|spim1_inst~O_SPI_MASTER_SCLK ;

assign hps_io_hps_io_spim1_inst_SS0 = \arm_a9_hps|hps_io|border|spim1_inst~O_SPI_MASTER_SS_0_N ;

assign hps_io_hps_io_uart0_inst_TX = \arm_a9_hps|hps_io|border|uart0_inst~uart_txd ;

assign memory_mem_a[0] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ;

assign memory_mem_a[1] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ;

assign memory_mem_a[2] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ;

assign memory_mem_a[3] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ;

assign memory_mem_a[4] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ;

assign memory_mem_a[5] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ;

assign memory_mem_a[6] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ;

assign memory_mem_a[7] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ;

assign memory_mem_a[8] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ;

assign memory_mem_a[9] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ;

assign memory_mem_a[10] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ;

assign memory_mem_a[11] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ;

assign memory_mem_a[12] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ;

assign memory_mem_a[13] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ;

assign memory_mem_a[14] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ;

assign memory_mem_ba[0] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ;

assign memory_mem_ba[1] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ;

assign memory_mem_ba[2] = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ;

assign memory_mem_cke = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ;

assign memory_mem_cs_n = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ;

assign memory_mem_ras_n = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ;

assign memory_mem_cas_n = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ;

assign memory_mem_we_n = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ;

assign memory_mem_reset_n = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ;

assign memory_mem_odt = \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ;

assign onchip_sram_s1_readdata[0] = \onchip_sram|the_altsyncram|auto_generated|q_a[0] ;

assign onchip_sram_s1_readdata[1] = \onchip_sram|the_altsyncram|auto_generated|q_a[1] ;

assign onchip_sram_s1_readdata[2] = \onchip_sram|the_altsyncram|auto_generated|q_a[2] ;

assign onchip_sram_s1_readdata[3] = \onchip_sram|the_altsyncram|auto_generated|q_a[3] ;

assign onchip_sram_s1_readdata[4] = \onchip_sram|the_altsyncram|auto_generated|q_a[4] ;

assign onchip_sram_s1_readdata[5] = \onchip_sram|the_altsyncram|auto_generated|q_a[5] ;

assign onchip_sram_s1_readdata[6] = \onchip_sram|the_altsyncram|auto_generated|q_a[6] ;

assign onchip_sram_s1_readdata[7] = \onchip_sram|the_altsyncram|auto_generated|q_a[7] ;

assign onchip_sram_s1_readdata[8] = \onchip_sram|the_altsyncram|auto_generated|q_a[8] ;

assign onchip_sram_s1_readdata[9] = \onchip_sram|the_altsyncram|auto_generated|q_a[9] ;

assign onchip_sram_s1_readdata[10] = \onchip_sram|the_altsyncram|auto_generated|q_a[10] ;

assign onchip_sram_s1_readdata[11] = \onchip_sram|the_altsyncram|auto_generated|q_a[11] ;

assign onchip_sram_s1_readdata[12] = \onchip_sram|the_altsyncram|auto_generated|q_a[12] ;

assign onchip_sram_s1_readdata[13] = \onchip_sram|the_altsyncram|auto_generated|q_a[13] ;

assign onchip_sram_s1_readdata[14] = \onchip_sram|the_altsyncram|auto_generated|q_a[14] ;

assign onchip_sram_s1_readdata[15] = \onchip_sram|the_altsyncram|auto_generated|q_a[15] ;

assign onchip_sram_s1_readdata[16] = \onchip_sram|the_altsyncram|auto_generated|q_a[16] ;

assign onchip_sram_s1_readdata[17] = \onchip_sram|the_altsyncram|auto_generated|q_a[17] ;

assign onchip_sram_s1_readdata[18] = \onchip_sram|the_altsyncram|auto_generated|q_a[18] ;

assign onchip_sram_s1_readdata[19] = \onchip_sram|the_altsyncram|auto_generated|q_a[19] ;

assign onchip_sram_s1_readdata[20] = \onchip_sram|the_altsyncram|auto_generated|q_a[20] ;

assign onchip_sram_s1_readdata[21] = \onchip_sram|the_altsyncram|auto_generated|q_a[21] ;

assign onchip_sram_s1_readdata[22] = \onchip_sram|the_altsyncram|auto_generated|q_a[22] ;

assign onchip_sram_s1_readdata[23] = \onchip_sram|the_altsyncram|auto_generated|q_a[23] ;

assign onchip_sram_s1_readdata[24] = \onchip_sram|the_altsyncram|auto_generated|q_a[24] ;

assign onchip_sram_s1_readdata[25] = \onchip_sram|the_altsyncram|auto_generated|q_a[25] ;

assign onchip_sram_s1_readdata[26] = \onchip_sram|the_altsyncram|auto_generated|q_a[26] ;

assign onchip_sram_s1_readdata[27] = \onchip_sram|the_altsyncram|auto_generated|q_a[27] ;

assign onchip_sram_s1_readdata[28] = \onchip_sram|the_altsyncram|auto_generated|q_a[28] ;

assign onchip_sram_s1_readdata[29] = \onchip_sram|the_altsyncram|auto_generated|q_a[29] ;

assign onchip_sram_s1_readdata[30] = \onchip_sram|the_altsyncram|auto_generated|q_a[30] ;

assign onchip_sram_s1_readdata[31] = \onchip_sram|the_altsyncram|auto_generated|q_a[31] ;

assign sdram_clk_clk = \system_pll|sys_pll|altera_pll_i|outclk_wire[1] ;

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[0] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[1] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_emac1_inst_MDIO),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[2] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[3] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO0),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO0[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[4] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[5] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO1),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO1[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[6] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[7] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO2),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO2[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[8] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[9] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_qspi_inst_IO3),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_qspi_inst_IO3[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[10] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[11] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_CMD),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_CMD[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[12] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[13] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D0),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D0[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[14] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[15] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D1),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D1[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[16] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[17] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D2),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D2[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[18] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[19] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_sdio_inst_D3),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_sdio_inst_D3[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[20] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[21] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D0),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D0[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[22] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[23] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D1),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D1[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[24] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[25] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D2),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D2[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[26] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[27] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D3),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D3[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[28] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[29] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D4),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D4[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[30] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[31] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D5),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D5[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[32] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[33] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D6),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D6[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[34] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[35] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_usb1_inst_D7),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_usb1_inst_D7[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~output (
	.i(!\arm_a9_hps|hps_io|border|intermediate[38] ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_i2c0_inst_SDA),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~output .open_drain_output = "true";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SDA[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~output (
	.i(!\arm_a9_hps|hps_io|border|intermediate[39] ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_i2c0_inst_SCL),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~output .open_drain_output = "true";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c0_inst_SCL[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~output (
	.i(!\arm_a9_hps|hps_io|border|intermediate[40] ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_i2c1_inst_SDA),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~output .open_drain_output = "true";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SDA[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~output (
	.i(!\arm_a9_hps|hps_io|border|intermediate[41] ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_i2c1_inst_SCL),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~output .open_drain_output = "true";
defparam \arm_a9_hps|hps_io|border|hps_io_i2c1_inst_SCL[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[42] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[43] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO09),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO09[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[44] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[45] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO35),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO35[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[46] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[47] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO40),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO40[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[48] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[49] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO41),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO41[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[50] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[51] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO48),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO48[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[52] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[53] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO53),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO53[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[54] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[55] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO54),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO54[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~output (
	.i(\arm_a9_hps|hps_io|border|intermediate[56] ),
	.oe(\arm_a9_hps|hps_io|border|intermediate[57] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_io_hps_io_gpio_inst_GPIO61),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~output .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~output .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_io_gpio_inst_GPIO61[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[0]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[1]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[2]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[3]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[4]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[5]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[6]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[7]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[8]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[9]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[10]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[11]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[12]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[13]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[14]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[15]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[16]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[17]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[18]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[19]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[20]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[21]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[22]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[23]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[24]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[25]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[26]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[27]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[28]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[29]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[30]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[31]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[0]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[1]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[2]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[3]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[0]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[1]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[2]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\arm_a9_hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[3]),
	.obar());
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \arm_a9_hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

endmodule

module Computer_System_altera_reset_controller (
	r_sync_rst1,
	r_early_rst1,
	merged_reset,
	clock_bridge_0_in_clk_clk)/* synthesis synthesis_greybox=0 */;
output 	r_sync_rst1;
output 	r_early_rst1;
input 	merged_reset;
input 	clock_bridge_0_in_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;
wire \always2~0_combout ;


Computer_System_altera_reset_synchronizer_4 alt_rst_req_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk(clock_bridge_0_in_clk_clk));

Computer_System_altera_reset_synchronizer_5 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.merged_reset(merged_reset),
	.clk(clock_bridge_0_in_clk_clk));

dffeas r_sync_rst(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas r_early_rst(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \altera_reset_synchronizer_int_chain[4]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~1 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~1 .extended_lut = "off";
defparam \r_sync_rst_chain~1 .lut_mask = 64'h1111111111111111;
defparam \r_sync_rst_chain~1 .shared_arith = "off";

dffeas \r_sync_rst_chain[2] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~0 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~0 .extended_lut = "off";
defparam \r_sync_rst_chain~0 .lut_mask = 64'h1111111111111111;
defparam \r_sync_rst_chain~0 .shared_arith = "off";

dffeas \r_sync_rst_chain[1] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!r_sync_rst1),
	.datab(!\altera_reset_synchronizer_int_chain[4]~q ),
	.datac(!\r_sync_rst_chain[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h7373737373737373;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always2~0 .shared_arith = "off";

endmodule

module Computer_System_altera_reset_controller_1 (
	h2f_rst_n_0,
	outclk_wire_0,
	locked_wire_0,
	r_early_rst1,
	r_sync_rst1,
	merged_reset)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
input 	outclk_wire_0;
input 	locked_wire_0;
output 	r_early_rst1;
output 	r_sync_rst1;
output 	merged_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \always2~0_combout ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;


Computer_System_altera_reset_synchronizer alt_rst_req_sync_uq1(
	.clk(outclk_wire_0),
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ));

Computer_System_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.clk(outclk_wire_0),
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.merged_reset(merged_reset));

dffeas r_early_rst(
	.clk(outclk_wire_0),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas r_sync_rst(
	.clk(outclk_wire_0),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

cyclonev_lcell_comb \merged_reset~0 (
	.dataa(!h2f_rst_n_0),
	.datab(!locked_wire_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(merged_reset),
	.sumout(),
	.cout(),
	.shareout());
defparam \merged_reset~0 .extended_lut = "off";
defparam \merged_reset~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \merged_reset~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(outclk_wire_0),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(outclk_wire_0),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(outclk_wire_0),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(outclk_wire_0),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~0 .extended_lut = "off";
defparam \r_sync_rst_chain~0 .lut_mask = 64'h1111111111111111;
defparam \r_sync_rst_chain~0 .shared_arith = "off";

dffeas \r_sync_rst_chain[2] (
	.clk(outclk_wire_0),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always2~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(outclk_wire_0),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \altera_reset_synchronizer_int_chain[4]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(outclk_wire_0),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~1 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~1 .extended_lut = "off";
defparam \r_sync_rst_chain~1 .lut_mask = 64'h1111111111111111;
defparam \r_sync_rst_chain~1 .shared_arith = "off";

dffeas \r_sync_rst_chain[1] (
	.clk(outclk_wire_0),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!r_sync_rst1),
	.datab(!\altera_reset_synchronizer_int_chain[4]~q ),
	.datac(!\r_sync_rst_chain[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h7373737373737373;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module Computer_System_altera_reset_synchronizer (
	clk,
	altera_reset_synchronizer_int_chain_out1)/* synthesis synthesis_greybox=0 */;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 64'h0000000000000000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module Computer_System_altera_reset_synchronizer_1 (
	clk,
	altera_reset_synchronizer_int_chain_out1,
	merged_reset)/* synthesis synthesis_greybox=0 */;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;
input 	merged_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module Computer_System_altera_reset_controller_2 (
	h2f_rst_n_0,
	outclk_wire_0,
	altera_reset_synchronizer_int_chain_out)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
input 	outclk_wire_0;
output 	altera_reset_synchronizer_int_chain_out;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altera_reset_synchronizer_3 alt_rst_sync_uq1(
	.h2f_rst_n_0(h2f_rst_n_0),
	.clk(outclk_wire_0),
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out));

endmodule

module Computer_System_altera_reset_synchronizer_3 (
	h2f_rst_n_0,
	clk,
	altera_reset_synchronizer_int_chain_out1)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
input 	clk;
output 	altera_reset_synchronizer_int_chain_out1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module Computer_System_altera_reset_synchronizer_4 (
	altera_reset_synchronizer_int_chain_out1,
	clk)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 64'h0000000000000000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module Computer_System_altera_reset_synchronizer_5 (
	altera_reset_synchronizer_int_chain_out1,
	merged_reset,
	clk)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	merged_reset;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module Computer_System_Computer_System_ARM_A9_HPS (
	h2f_rst_n_0,
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	h2f_ARVALID_0,
	h2f_AWVALID_0,
	h2f_BREADY_0,
	h2f_RREADY_0,
	h2f_WLAST_0,
	h2f_WVALID_0,
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARADDR_4,
	h2f_ARADDR_5,
	h2f_ARADDR_6,
	h2f_ARADDR_7,
	h2f_ARADDR_8,
	h2f_ARADDR_9,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARLEN_0,
	h2f_ARLEN_1,
	h2f_ARLEN_2,
	h2f_ARLEN_3,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWADDR_0,
	h2f_AWADDR_1,
	h2f_AWADDR_2,
	h2f_AWADDR_3,
	h2f_AWADDR_4,
	h2f_AWADDR_5,
	h2f_AWADDR_6,
	h2f_AWADDR_7,
	h2f_AWADDR_8,
	h2f_AWADDR_9,
	h2f_AWADDR_10,
	h2f_AWADDR_11,
	h2f_AWADDR_12,
	h2f_AWADDR_13,
	h2f_AWADDR_14,
	h2f_AWADDR_15,
	h2f_AWADDR_16,
	h2f_AWADDR_17,
	h2f_AWADDR_18,
	h2f_AWADDR_19,
	h2f_AWADDR_20,
	h2f_AWADDR_21,
	h2f_AWADDR_22,
	h2f_AWADDR_23,
	h2f_AWADDR_24,
	h2f_AWADDR_25,
	h2f_AWADDR_26,
	h2f_AWADDR_27,
	h2f_AWBURST_0,
	h2f_AWBURST_1,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWLEN_0,
	h2f_AWLEN_1,
	h2f_AWLEN_2,
	h2f_AWLEN_3,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WDATA_1,
	h2f_WDATA_2,
	h2f_WDATA_3,
	h2f_WDATA_4,
	h2f_WDATA_5,
	h2f_WDATA_6,
	h2f_WDATA_7,
	h2f_WDATA_8,
	h2f_WDATA_9,
	h2f_WDATA_10,
	h2f_WDATA_11,
	h2f_WDATA_12,
	h2f_WDATA_13,
	h2f_WDATA_14,
	h2f_WDATA_15,
	h2f_WDATA_16,
	h2f_WDATA_17,
	h2f_WDATA_18,
	h2f_WDATA_19,
	h2f_WDATA_20,
	h2f_WDATA_21,
	h2f_WDATA_22,
	h2f_WDATA_23,
	h2f_WDATA_24,
	h2f_WDATA_25,
	h2f_WDATA_26,
	h2f_WDATA_27,
	h2f_WDATA_28,
	h2f_WDATA_29,
	h2f_WDATA_30,
	h2f_WDATA_31,
	h2f_WDATA_32,
	h2f_WDATA_33,
	h2f_WDATA_34,
	h2f_WDATA_35,
	h2f_WDATA_36,
	h2f_WDATA_37,
	h2f_WDATA_38,
	h2f_WDATA_39,
	h2f_WDATA_40,
	h2f_WDATA_41,
	h2f_WDATA_42,
	h2f_WDATA_43,
	h2f_WDATA_44,
	h2f_WDATA_45,
	h2f_WDATA_46,
	h2f_WDATA_47,
	h2f_WDATA_48,
	h2f_WDATA_49,
	h2f_WDATA_50,
	h2f_WDATA_51,
	h2f_WDATA_52,
	h2f_WDATA_53,
	h2f_WDATA_54,
	h2f_WDATA_55,
	h2f_WDATA_56,
	h2f_WDATA_57,
	h2f_WDATA_58,
	h2f_WDATA_59,
	h2f_WDATA_60,
	h2f_WDATA_61,
	h2f_WDATA_62,
	h2f_WDATA_63,
	h2f_WDATA_64,
	h2f_WDATA_65,
	h2f_WDATA_66,
	h2f_WDATA_67,
	h2f_WDATA_68,
	h2f_WDATA_69,
	h2f_WDATA_70,
	h2f_WDATA_71,
	h2f_WDATA_72,
	h2f_WDATA_73,
	h2f_WDATA_74,
	h2f_WDATA_75,
	h2f_WDATA_76,
	h2f_WDATA_77,
	h2f_WDATA_78,
	h2f_WDATA_79,
	h2f_WDATA_80,
	h2f_WDATA_81,
	h2f_WDATA_82,
	h2f_WDATA_83,
	h2f_WDATA_84,
	h2f_WDATA_85,
	h2f_WDATA_86,
	h2f_WDATA_87,
	h2f_WDATA_88,
	h2f_WDATA_89,
	h2f_WDATA_90,
	h2f_WDATA_91,
	h2f_WDATA_92,
	h2f_WDATA_93,
	h2f_WDATA_94,
	h2f_WDATA_95,
	h2f_WDATA_96,
	h2f_WDATA_97,
	h2f_WDATA_98,
	h2f_WDATA_99,
	h2f_WDATA_100,
	h2f_WDATA_101,
	h2f_WDATA_102,
	h2f_WDATA_103,
	h2f_WDATA_104,
	h2f_WDATA_105,
	h2f_WDATA_106,
	h2f_WDATA_107,
	h2f_WDATA_108,
	h2f_WDATA_109,
	h2f_WDATA_110,
	h2f_WDATA_111,
	h2f_WDATA_112,
	h2f_WDATA_113,
	h2f_WDATA_114,
	h2f_WDATA_115,
	h2f_WDATA_116,
	h2f_WDATA_117,
	h2f_WDATA_118,
	h2f_WDATA_119,
	h2f_WDATA_120,
	h2f_WDATA_121,
	h2f_WDATA_122,
	h2f_WDATA_123,
	h2f_WDATA_124,
	h2f_WDATA_125,
	h2f_WDATA_126,
	h2f_WDATA_127,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	h2f_WSTRB_4,
	h2f_WSTRB_5,
	h2f_WSTRB_6,
	h2f_WSTRB_7,
	h2f_WSTRB_8,
	h2f_WSTRB_9,
	h2f_WSTRB_10,
	h2f_WSTRB_11,
	h2f_WSTRB_12,
	h2f_WSTRB_13,
	h2f_WSTRB_14,
	h2f_WSTRB_15,
	outclk_wire_0,
	sink1_ready,
	awready,
	src0_valid,
	source_endofpacket,
	src1_valid,
	wready,
	mem_88_0,
	mem_89_0,
	mem_90_0,
	mem_91_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	sink1_ready1,
	awready1,
	WideOr1,
	src_payload_0,
	WideOr11,
	wready1,
	src_data_209,
	src_data_210,
	src_data_211,
	src_data_212,
	src_data_213,
	src_data_214,
	src_data_215,
	src_data_216,
	src_data_217,
	src_data_218,
	src_data_219,
	src_data_220,
	src_data_0,
	src_payload,
	src_data_2,
	src_data_3,
	src_payload1,
	src_data_5,
	src_payload2,
	src_data_7,
	src_payload3,
	src_data_9,
	src_data_10,
	src_data_11,
	src_data_12,
	src_payload4,
	src_data_14,
	src_data_15,
	src_data_16,
	src_payload5,
	src_data_18,
	src_data_19,
	src_payload6,
	src_data_21,
	src_payload7,
	src_data_23,
	src_payload8,
	src_data_25,
	src_data_26,
	src_data_27,
	src_data_28,
	src_payload9,
	src_data_30,
	src_data_31,
	src_data_32,
	src_payload10,
	src_data_34,
	src_data_35,
	src_payload11,
	src_data_37,
	src_payload12,
	src_data_39,
	src_payload13,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_payload14,
	src_data_46,
	src_data_47,
	src_data_48,
	src_payload15,
	src_data_50,
	src_data_51,
	src_payload16,
	src_data_53,
	src_payload17,
	src_data_55,
	src_payload18,
	src_data_57,
	src_data_58,
	src_data_59,
	src_data_60,
	src_payload19,
	src_data_62,
	src_data_63,
	src_data_64,
	src_payload20,
	src_data_66,
	src_data_67,
	src_payload21,
	src_data_69,
	src_payload22,
	src_data_71,
	src_payload23,
	src_data_73,
	src_data_74,
	src_data_75,
	src_data_76,
	src_payload24,
	src_data_78,
	src_data_79,
	src_data_80,
	src_payload25,
	src_data_82,
	src_data_83,
	src_payload26,
	src_data_85,
	src_payload27,
	src_data_87,
	src_payload28,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_payload29,
	src_data_94,
	src_data_95,
	src_data_96,
	src_payload30,
	src_data_98,
	src_data_99,
	src_payload31,
	src_data_101,
	src_payload32,
	src_data_103,
	src_payload33,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_payload34,
	src_data_110,
	src_data_111,
	src_data_112,
	src_payload35,
	src_data_114,
	src_data_115,
	src_payload36,
	src_data_117,
	src_payload37,
	src_data_119,
	src_payload38,
	src_data_121,
	src_data_122,
	src_data_123,
	src_data_124,
	src_payload39,
	src_data_126,
	src_data_127,
	src_data_2091,
	src_data_2101,
	src_data_2111,
	src_data_2121,
	src_data_2131,
	src_data_2141,
	src_data_2151,
	src_data_2161,
	src_data_2171,
	src_data_2181,
	src_data_2191,
	src_data_2201,
	emac1_inst,
	emac1_inst1,
	intermediate_0,
	intermediate_1,
	emac1_inst2,
	emac1_inst3,
	emac1_inst4,
	emac1_inst5,
	emac1_inst6,
	qspi_inst,
	intermediate_2,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_3,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	qspi_inst1,
	sdio_inst,
	intermediate_10,
	intermediate_11,
	intermediate_12,
	intermediate_14,
	intermediate_16,
	intermediate_18,
	intermediate_13,
	intermediate_15,
	intermediate_17,
	intermediate_19,
	usb1_inst,
	intermediate_20,
	intermediate_22,
	intermediate_24,
	intermediate_26,
	intermediate_28,
	intermediate_30,
	intermediate_32,
	intermediate_34,
	intermediate_21,
	intermediate_23,
	intermediate_25,
	intermediate_27,
	intermediate_29,
	intermediate_31,
	intermediate_33,
	intermediate_35,
	spim1_inst,
	spim1_inst1,
	intermediate_36,
	intermediate_37,
	uart0_inst,
	intermediate_39,
	intermediate_38,
	intermediate_41,
	intermediate_40,
	intermediate_42,
	intermediate_43,
	intermediate_44,
	intermediate_46,
	intermediate_48,
	intermediate_50,
	intermediate_52,
	intermediate_54,
	intermediate_45,
	intermediate_47,
	intermediate_49,
	intermediate_51,
	intermediate_53,
	intermediate_55,
	intermediate_56,
	intermediate_57,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_qspi_inst_IO0_0,
	hps_io_qspi_inst_IO1_0,
	hps_io_qspi_inst_IO2_0,
	hps_io_qspi_inst_IO3_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_io_usb1_inst_D0_0,
	hps_io_usb1_inst_D1_0,
	hps_io_usb1_inst_D2_0,
	hps_io_usb1_inst_D3_0,
	hps_io_usb1_inst_D4_0,
	hps_io_usb1_inst_D5_0,
	hps_io_usb1_inst_D6_0,
	hps_io_usb1_inst_D7_0,
	hps_io_i2c0_inst_SDA_0,
	hps_io_i2c0_inst_SCL_0,
	hps_io_i2c1_inst_SDA_0,
	hps_io_i2c1_inst_SCL_0,
	hps_io_gpio_inst_GPIO09_0,
	hps_io_gpio_inst_GPIO35_0,
	hps_io_gpio_inst_GPIO40_0,
	hps_io_gpio_inst_GPIO41_0,
	hps_io_gpio_inst_GPIO48_0,
	hps_io_gpio_inst_GPIO53_0,
	hps_io_gpio_inst_GPIO54_0,
	hps_io_gpio_inst_GPIO61_0,
	hps_io_hps_io_emac1_inst_RXD0,
	hps_io_hps_io_emac1_inst_RXD1,
	hps_io_hps_io_emac1_inst_RXD2,
	hps_io_hps_io_emac1_inst_RXD3,
	hps_io_hps_io_emac1_inst_RX_CLK,
	hps_io_hps_io_emac1_inst_RX_CTL,
	hps_io_hps_io_spim1_inst_MISO,
	hps_io_hps_io_uart0_inst_RX,
	hps_io_hps_io_usb1_inst_CLK,
	hps_io_hps_io_usb1_inst_DIR,
	hps_io_hps_io_usb1_inst_NXT,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	h2f_rst_n_0;
output 	h2f_lw_ARVALID_0;
output 	h2f_lw_AWVALID_0;
output 	h2f_lw_BREADY_0;
output 	h2f_lw_RREADY_0;
output 	h2f_lw_WLAST_0;
output 	h2f_lw_WVALID_0;
output 	h2f_lw_ARADDR_0;
output 	h2f_lw_ARADDR_1;
output 	h2f_lw_ARADDR_2;
output 	h2f_lw_ARADDR_3;
output 	h2f_lw_ARADDR_4;
output 	h2f_lw_ARBURST_0;
output 	h2f_lw_ARBURST_1;
output 	h2f_lw_ARID_0;
output 	h2f_lw_ARID_1;
output 	h2f_lw_ARID_2;
output 	h2f_lw_ARID_3;
output 	h2f_lw_ARID_4;
output 	h2f_lw_ARID_5;
output 	h2f_lw_ARID_6;
output 	h2f_lw_ARID_7;
output 	h2f_lw_ARID_8;
output 	h2f_lw_ARID_9;
output 	h2f_lw_ARID_10;
output 	h2f_lw_ARID_11;
output 	h2f_lw_ARLEN_0;
output 	h2f_lw_ARLEN_1;
output 	h2f_lw_ARLEN_2;
output 	h2f_lw_ARLEN_3;
output 	h2f_lw_ARSIZE_0;
output 	h2f_lw_ARSIZE_1;
output 	h2f_lw_ARSIZE_2;
output 	h2f_lw_AWADDR_0;
output 	h2f_lw_AWADDR_1;
output 	h2f_lw_AWADDR_2;
output 	h2f_lw_AWADDR_3;
output 	h2f_lw_AWADDR_4;
output 	h2f_lw_AWBURST_0;
output 	h2f_lw_AWBURST_1;
output 	h2f_lw_AWID_0;
output 	h2f_lw_AWID_1;
output 	h2f_lw_AWID_2;
output 	h2f_lw_AWID_3;
output 	h2f_lw_AWID_4;
output 	h2f_lw_AWID_5;
output 	h2f_lw_AWID_6;
output 	h2f_lw_AWID_7;
output 	h2f_lw_AWID_8;
output 	h2f_lw_AWID_9;
output 	h2f_lw_AWID_10;
output 	h2f_lw_AWID_11;
output 	h2f_lw_AWLEN_0;
output 	h2f_lw_AWLEN_1;
output 	h2f_lw_AWLEN_2;
output 	h2f_lw_AWLEN_3;
output 	h2f_lw_AWSIZE_0;
output 	h2f_lw_AWSIZE_1;
output 	h2f_lw_AWSIZE_2;
output 	h2f_lw_WDATA_0;
output 	h2f_lw_WDATA_1;
output 	h2f_lw_WDATA_2;
output 	h2f_lw_WDATA_3;
output 	h2f_lw_WDATA_4;
output 	h2f_lw_WDATA_5;
output 	h2f_lw_WDATA_6;
output 	h2f_lw_WDATA_7;
output 	h2f_lw_WDATA_8;
output 	h2f_lw_WDATA_9;
output 	h2f_lw_WDATA_10;
output 	h2f_lw_WDATA_11;
output 	h2f_lw_WDATA_12;
output 	h2f_lw_WDATA_13;
output 	h2f_lw_WDATA_14;
output 	h2f_lw_WDATA_15;
output 	h2f_lw_WDATA_16;
output 	h2f_lw_WDATA_17;
output 	h2f_lw_WDATA_18;
output 	h2f_lw_WDATA_19;
output 	h2f_lw_WDATA_20;
output 	h2f_lw_WDATA_21;
output 	h2f_lw_WDATA_22;
output 	h2f_lw_WDATA_23;
output 	h2f_lw_WDATA_24;
output 	h2f_lw_WDATA_25;
output 	h2f_lw_WDATA_26;
output 	h2f_lw_WDATA_27;
output 	h2f_lw_WDATA_28;
output 	h2f_lw_WDATA_29;
output 	h2f_lw_WDATA_30;
output 	h2f_lw_WDATA_31;
output 	h2f_lw_WSTRB_0;
output 	h2f_lw_WSTRB_1;
output 	h2f_lw_WSTRB_2;
output 	h2f_lw_WSTRB_3;
output 	h2f_ARVALID_0;
output 	h2f_AWVALID_0;
output 	h2f_BREADY_0;
output 	h2f_RREADY_0;
output 	h2f_WLAST_0;
output 	h2f_WVALID_0;
output 	h2f_ARADDR_0;
output 	h2f_ARADDR_1;
output 	h2f_ARADDR_2;
output 	h2f_ARADDR_3;
output 	h2f_ARADDR_4;
output 	h2f_ARADDR_5;
output 	h2f_ARADDR_6;
output 	h2f_ARADDR_7;
output 	h2f_ARADDR_8;
output 	h2f_ARADDR_9;
output 	h2f_ARBURST_0;
output 	h2f_ARBURST_1;
output 	h2f_ARID_0;
output 	h2f_ARID_1;
output 	h2f_ARID_2;
output 	h2f_ARID_3;
output 	h2f_ARID_4;
output 	h2f_ARID_5;
output 	h2f_ARID_6;
output 	h2f_ARID_7;
output 	h2f_ARID_8;
output 	h2f_ARID_9;
output 	h2f_ARID_10;
output 	h2f_ARID_11;
output 	h2f_ARLEN_0;
output 	h2f_ARLEN_1;
output 	h2f_ARLEN_2;
output 	h2f_ARLEN_3;
output 	h2f_ARSIZE_0;
output 	h2f_ARSIZE_1;
output 	h2f_ARSIZE_2;
output 	h2f_AWADDR_0;
output 	h2f_AWADDR_1;
output 	h2f_AWADDR_2;
output 	h2f_AWADDR_3;
output 	h2f_AWADDR_4;
output 	h2f_AWADDR_5;
output 	h2f_AWADDR_6;
output 	h2f_AWADDR_7;
output 	h2f_AWADDR_8;
output 	h2f_AWADDR_9;
output 	h2f_AWADDR_10;
output 	h2f_AWADDR_11;
output 	h2f_AWADDR_12;
output 	h2f_AWADDR_13;
output 	h2f_AWADDR_14;
output 	h2f_AWADDR_15;
output 	h2f_AWADDR_16;
output 	h2f_AWADDR_17;
output 	h2f_AWADDR_18;
output 	h2f_AWADDR_19;
output 	h2f_AWADDR_20;
output 	h2f_AWADDR_21;
output 	h2f_AWADDR_22;
output 	h2f_AWADDR_23;
output 	h2f_AWADDR_24;
output 	h2f_AWADDR_25;
output 	h2f_AWADDR_26;
output 	h2f_AWADDR_27;
output 	h2f_AWBURST_0;
output 	h2f_AWBURST_1;
output 	h2f_AWID_0;
output 	h2f_AWID_1;
output 	h2f_AWID_2;
output 	h2f_AWID_3;
output 	h2f_AWID_4;
output 	h2f_AWID_5;
output 	h2f_AWID_6;
output 	h2f_AWID_7;
output 	h2f_AWID_8;
output 	h2f_AWID_9;
output 	h2f_AWID_10;
output 	h2f_AWID_11;
output 	h2f_AWLEN_0;
output 	h2f_AWLEN_1;
output 	h2f_AWLEN_2;
output 	h2f_AWLEN_3;
output 	h2f_AWSIZE_0;
output 	h2f_AWSIZE_1;
output 	h2f_AWSIZE_2;
output 	h2f_WDATA_0;
output 	h2f_WDATA_1;
output 	h2f_WDATA_2;
output 	h2f_WDATA_3;
output 	h2f_WDATA_4;
output 	h2f_WDATA_5;
output 	h2f_WDATA_6;
output 	h2f_WDATA_7;
output 	h2f_WDATA_8;
output 	h2f_WDATA_9;
output 	h2f_WDATA_10;
output 	h2f_WDATA_11;
output 	h2f_WDATA_12;
output 	h2f_WDATA_13;
output 	h2f_WDATA_14;
output 	h2f_WDATA_15;
output 	h2f_WDATA_16;
output 	h2f_WDATA_17;
output 	h2f_WDATA_18;
output 	h2f_WDATA_19;
output 	h2f_WDATA_20;
output 	h2f_WDATA_21;
output 	h2f_WDATA_22;
output 	h2f_WDATA_23;
output 	h2f_WDATA_24;
output 	h2f_WDATA_25;
output 	h2f_WDATA_26;
output 	h2f_WDATA_27;
output 	h2f_WDATA_28;
output 	h2f_WDATA_29;
output 	h2f_WDATA_30;
output 	h2f_WDATA_31;
output 	h2f_WDATA_32;
output 	h2f_WDATA_33;
output 	h2f_WDATA_34;
output 	h2f_WDATA_35;
output 	h2f_WDATA_36;
output 	h2f_WDATA_37;
output 	h2f_WDATA_38;
output 	h2f_WDATA_39;
output 	h2f_WDATA_40;
output 	h2f_WDATA_41;
output 	h2f_WDATA_42;
output 	h2f_WDATA_43;
output 	h2f_WDATA_44;
output 	h2f_WDATA_45;
output 	h2f_WDATA_46;
output 	h2f_WDATA_47;
output 	h2f_WDATA_48;
output 	h2f_WDATA_49;
output 	h2f_WDATA_50;
output 	h2f_WDATA_51;
output 	h2f_WDATA_52;
output 	h2f_WDATA_53;
output 	h2f_WDATA_54;
output 	h2f_WDATA_55;
output 	h2f_WDATA_56;
output 	h2f_WDATA_57;
output 	h2f_WDATA_58;
output 	h2f_WDATA_59;
output 	h2f_WDATA_60;
output 	h2f_WDATA_61;
output 	h2f_WDATA_62;
output 	h2f_WDATA_63;
output 	h2f_WDATA_64;
output 	h2f_WDATA_65;
output 	h2f_WDATA_66;
output 	h2f_WDATA_67;
output 	h2f_WDATA_68;
output 	h2f_WDATA_69;
output 	h2f_WDATA_70;
output 	h2f_WDATA_71;
output 	h2f_WDATA_72;
output 	h2f_WDATA_73;
output 	h2f_WDATA_74;
output 	h2f_WDATA_75;
output 	h2f_WDATA_76;
output 	h2f_WDATA_77;
output 	h2f_WDATA_78;
output 	h2f_WDATA_79;
output 	h2f_WDATA_80;
output 	h2f_WDATA_81;
output 	h2f_WDATA_82;
output 	h2f_WDATA_83;
output 	h2f_WDATA_84;
output 	h2f_WDATA_85;
output 	h2f_WDATA_86;
output 	h2f_WDATA_87;
output 	h2f_WDATA_88;
output 	h2f_WDATA_89;
output 	h2f_WDATA_90;
output 	h2f_WDATA_91;
output 	h2f_WDATA_92;
output 	h2f_WDATA_93;
output 	h2f_WDATA_94;
output 	h2f_WDATA_95;
output 	h2f_WDATA_96;
output 	h2f_WDATA_97;
output 	h2f_WDATA_98;
output 	h2f_WDATA_99;
output 	h2f_WDATA_100;
output 	h2f_WDATA_101;
output 	h2f_WDATA_102;
output 	h2f_WDATA_103;
output 	h2f_WDATA_104;
output 	h2f_WDATA_105;
output 	h2f_WDATA_106;
output 	h2f_WDATA_107;
output 	h2f_WDATA_108;
output 	h2f_WDATA_109;
output 	h2f_WDATA_110;
output 	h2f_WDATA_111;
output 	h2f_WDATA_112;
output 	h2f_WDATA_113;
output 	h2f_WDATA_114;
output 	h2f_WDATA_115;
output 	h2f_WDATA_116;
output 	h2f_WDATA_117;
output 	h2f_WDATA_118;
output 	h2f_WDATA_119;
output 	h2f_WDATA_120;
output 	h2f_WDATA_121;
output 	h2f_WDATA_122;
output 	h2f_WDATA_123;
output 	h2f_WDATA_124;
output 	h2f_WDATA_125;
output 	h2f_WDATA_126;
output 	h2f_WDATA_127;
output 	h2f_WSTRB_0;
output 	h2f_WSTRB_1;
output 	h2f_WSTRB_2;
output 	h2f_WSTRB_3;
output 	h2f_WSTRB_4;
output 	h2f_WSTRB_5;
output 	h2f_WSTRB_6;
output 	h2f_WSTRB_7;
output 	h2f_WSTRB_8;
output 	h2f_WSTRB_9;
output 	h2f_WSTRB_10;
output 	h2f_WSTRB_11;
output 	h2f_WSTRB_12;
output 	h2f_WSTRB_13;
output 	h2f_WSTRB_14;
output 	h2f_WSTRB_15;
input 	outclk_wire_0;
input 	sink1_ready;
input 	awready;
input 	src0_valid;
input 	source_endofpacket;
input 	src1_valid;
input 	wready;
input 	mem_88_0;
input 	mem_89_0;
input 	mem_90_0;
input 	mem_91_0;
input 	mem_92_0;
input 	mem_93_0;
input 	mem_94_0;
input 	mem_95_0;
input 	mem_96_0;
input 	mem_97_0;
input 	mem_98_0;
input 	mem_99_0;
input 	out_data_0;
input 	out_data_1;
input 	out_data_2;
input 	out_data_3;
input 	out_data_4;
input 	out_data_5;
input 	out_data_6;
input 	out_data_7;
input 	sink1_ready1;
input 	awready1;
input 	WideOr1;
input 	src_payload_0;
input 	WideOr11;
input 	wready1;
input 	src_data_209;
input 	src_data_210;
input 	src_data_211;
input 	src_data_212;
input 	src_data_213;
input 	src_data_214;
input 	src_data_215;
input 	src_data_216;
input 	src_data_217;
input 	src_data_218;
input 	src_data_219;
input 	src_data_220;
input 	src_data_0;
input 	src_payload;
input 	src_data_2;
input 	src_data_3;
input 	src_payload1;
input 	src_data_5;
input 	src_payload2;
input 	src_data_7;
input 	src_payload3;
input 	src_data_9;
input 	src_data_10;
input 	src_data_11;
input 	src_data_12;
input 	src_payload4;
input 	src_data_14;
input 	src_data_15;
input 	src_data_16;
input 	src_payload5;
input 	src_data_18;
input 	src_data_19;
input 	src_payload6;
input 	src_data_21;
input 	src_payload7;
input 	src_data_23;
input 	src_payload8;
input 	src_data_25;
input 	src_data_26;
input 	src_data_27;
input 	src_data_28;
input 	src_payload9;
input 	src_data_30;
input 	src_data_31;
input 	src_data_32;
input 	src_payload10;
input 	src_data_34;
input 	src_data_35;
input 	src_payload11;
input 	src_data_37;
input 	src_payload12;
input 	src_data_39;
input 	src_payload13;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_payload14;
input 	src_data_46;
input 	src_data_47;
input 	src_data_48;
input 	src_payload15;
input 	src_data_50;
input 	src_data_51;
input 	src_payload16;
input 	src_data_53;
input 	src_payload17;
input 	src_data_55;
input 	src_payload18;
input 	src_data_57;
input 	src_data_58;
input 	src_data_59;
input 	src_data_60;
input 	src_payload19;
input 	src_data_62;
input 	src_data_63;
input 	src_data_64;
input 	src_payload20;
input 	src_data_66;
input 	src_data_67;
input 	src_payload21;
input 	src_data_69;
input 	src_payload22;
input 	src_data_71;
input 	src_payload23;
input 	src_data_73;
input 	src_data_74;
input 	src_data_75;
input 	src_data_76;
input 	src_payload24;
input 	src_data_78;
input 	src_data_79;
input 	src_data_80;
input 	src_payload25;
input 	src_data_82;
input 	src_data_83;
input 	src_payload26;
input 	src_data_85;
input 	src_payload27;
input 	src_data_87;
input 	src_payload28;
input 	src_data_89;
input 	src_data_90;
input 	src_data_91;
input 	src_data_92;
input 	src_payload29;
input 	src_data_94;
input 	src_data_95;
input 	src_data_96;
input 	src_payload30;
input 	src_data_98;
input 	src_data_99;
input 	src_payload31;
input 	src_data_101;
input 	src_payload32;
input 	src_data_103;
input 	src_payload33;
input 	src_data_105;
input 	src_data_106;
input 	src_data_107;
input 	src_data_108;
input 	src_payload34;
input 	src_data_110;
input 	src_data_111;
input 	src_data_112;
input 	src_payload35;
input 	src_data_114;
input 	src_data_115;
input 	src_payload36;
input 	src_data_117;
input 	src_payload37;
input 	src_data_119;
input 	src_payload38;
input 	src_data_121;
input 	src_data_122;
input 	src_data_123;
input 	src_data_124;
input 	src_payload39;
input 	src_data_126;
input 	src_data_127;
input 	src_data_2091;
input 	src_data_2101;
input 	src_data_2111;
input 	src_data_2121;
input 	src_data_2131;
input 	src_data_2141;
input 	src_data_2151;
input 	src_data_2161;
input 	src_data_2171;
input 	src_data_2181;
input 	src_data_2191;
input 	src_data_2201;
output 	emac1_inst;
output 	emac1_inst1;
output 	intermediate_0;
output 	intermediate_1;
output 	emac1_inst2;
output 	emac1_inst3;
output 	emac1_inst4;
output 	emac1_inst5;
output 	emac1_inst6;
output 	qspi_inst;
output 	intermediate_2;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_3;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	qspi_inst1;
output 	sdio_inst;
output 	intermediate_10;
output 	intermediate_11;
output 	intermediate_12;
output 	intermediate_14;
output 	intermediate_16;
output 	intermediate_18;
output 	intermediate_13;
output 	intermediate_15;
output 	intermediate_17;
output 	intermediate_19;
output 	usb1_inst;
output 	intermediate_20;
output 	intermediate_22;
output 	intermediate_24;
output 	intermediate_26;
output 	intermediate_28;
output 	intermediate_30;
output 	intermediate_32;
output 	intermediate_34;
output 	intermediate_21;
output 	intermediate_23;
output 	intermediate_25;
output 	intermediate_27;
output 	intermediate_29;
output 	intermediate_31;
output 	intermediate_33;
output 	intermediate_35;
output 	spim1_inst;
output 	spim1_inst1;
output 	intermediate_36;
output 	intermediate_37;
output 	uart0_inst;
output 	intermediate_39;
output 	intermediate_38;
output 	intermediate_41;
output 	intermediate_40;
output 	intermediate_42;
output 	intermediate_43;
output 	intermediate_44;
output 	intermediate_46;
output 	intermediate_48;
output 	intermediate_50;
output 	intermediate_52;
output 	intermediate_54;
output 	intermediate_45;
output 	intermediate_47;
output 	intermediate_49;
output 	intermediate_51;
output 	intermediate_53;
output 	intermediate_55;
output 	intermediate_56;
output 	intermediate_57;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_qspi_inst_IO0_0;
input 	hps_io_qspi_inst_IO1_0;
input 	hps_io_qspi_inst_IO2_0;
input 	hps_io_qspi_inst_IO3_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_io_usb1_inst_D0_0;
input 	hps_io_usb1_inst_D1_0;
input 	hps_io_usb1_inst_D2_0;
input 	hps_io_usb1_inst_D3_0;
input 	hps_io_usb1_inst_D4_0;
input 	hps_io_usb1_inst_D5_0;
input 	hps_io_usb1_inst_D6_0;
input 	hps_io_usb1_inst_D7_0;
input 	hps_io_i2c0_inst_SDA_0;
input 	hps_io_i2c0_inst_SCL_0;
input 	hps_io_i2c1_inst_SDA_0;
input 	hps_io_i2c1_inst_SCL_0;
input 	hps_io_gpio_inst_GPIO09_0;
input 	hps_io_gpio_inst_GPIO35_0;
input 	hps_io_gpio_inst_GPIO40_0;
input 	hps_io_gpio_inst_GPIO41_0;
input 	hps_io_gpio_inst_GPIO48_0;
input 	hps_io_gpio_inst_GPIO53_0;
input 	hps_io_gpio_inst_GPIO54_0;
input 	hps_io_gpio_inst_GPIO61_0;
input 	hps_io_hps_io_emac1_inst_RXD0;
input 	hps_io_hps_io_emac1_inst_RXD1;
input 	hps_io_hps_io_emac1_inst_RXD2;
input 	hps_io_hps_io_emac1_inst_RXD3;
input 	hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_io_hps_io_emac1_inst_RX_CTL;
input 	hps_io_hps_io_spim1_inst_MISO;
input 	hps_io_hps_io_uart0_inst_RX;
input 	hps_io_hps_io_usb1_inst_CLK;
input 	hps_io_hps_io_usb1_inst_DIR;
input 	hps_io_hps_io_usb1_inst_NXT;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_Computer_System_ARM_A9_HPS_hps_io hps_io(
	.emac1_inst(emac1_inst),
	.emac1_inst1(emac1_inst1),
	.intermediate_0(intermediate_0),
	.intermediate_1(intermediate_1),
	.emac1_inst2(emac1_inst2),
	.emac1_inst3(emac1_inst3),
	.emac1_inst4(emac1_inst4),
	.emac1_inst5(emac1_inst5),
	.emac1_inst6(emac1_inst6),
	.qspi_inst(qspi_inst),
	.intermediate_2(intermediate_2),
	.intermediate_4(intermediate_4),
	.intermediate_6(intermediate_6),
	.intermediate_8(intermediate_8),
	.intermediate_3(intermediate_3),
	.intermediate_5(intermediate_5),
	.intermediate_7(intermediate_7),
	.intermediate_9(intermediate_9),
	.qspi_inst1(qspi_inst1),
	.sdio_inst(sdio_inst),
	.intermediate_10(intermediate_10),
	.intermediate_11(intermediate_11),
	.intermediate_12(intermediate_12),
	.intermediate_14(intermediate_14),
	.intermediate_16(intermediate_16),
	.intermediate_18(intermediate_18),
	.intermediate_13(intermediate_13),
	.intermediate_15(intermediate_15),
	.intermediate_17(intermediate_17),
	.intermediate_19(intermediate_19),
	.usb1_inst(usb1_inst),
	.intermediate_20(intermediate_20),
	.intermediate_22(intermediate_22),
	.intermediate_24(intermediate_24),
	.intermediate_26(intermediate_26),
	.intermediate_28(intermediate_28),
	.intermediate_30(intermediate_30),
	.intermediate_32(intermediate_32),
	.intermediate_34(intermediate_34),
	.intermediate_21(intermediate_21),
	.intermediate_23(intermediate_23),
	.intermediate_25(intermediate_25),
	.intermediate_27(intermediate_27),
	.intermediate_29(intermediate_29),
	.intermediate_31(intermediate_31),
	.intermediate_33(intermediate_33),
	.intermediate_35(intermediate_35),
	.spim1_inst(spim1_inst),
	.spim1_inst1(spim1_inst1),
	.intermediate_36(intermediate_36),
	.intermediate_37(intermediate_37),
	.uart0_inst(uart0_inst),
	.intermediate_39(intermediate_39),
	.intermediate_38(intermediate_38),
	.intermediate_41(intermediate_41),
	.intermediate_40(intermediate_40),
	.intermediate_42(intermediate_42),
	.intermediate_43(intermediate_43),
	.intermediate_44(intermediate_44),
	.intermediate_46(intermediate_46),
	.intermediate_48(intermediate_48),
	.intermediate_50(intermediate_50),
	.intermediate_52(intermediate_52),
	.intermediate_54(intermediate_54),
	.intermediate_45(intermediate_45),
	.intermediate_47(intermediate_47),
	.intermediate_49(intermediate_49),
	.intermediate_51(intermediate_51),
	.intermediate_53(intermediate_53),
	.intermediate_55(intermediate_55),
	.intermediate_56(intermediate_56),
	.intermediate_57(intermediate_57),
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.hps_io_emac1_inst_MDIO_0(hps_io_emac1_inst_MDIO_0),
	.hps_io_qspi_inst_IO0_0(hps_io_qspi_inst_IO0_0),
	.hps_io_qspi_inst_IO1_0(hps_io_qspi_inst_IO1_0),
	.hps_io_qspi_inst_IO2_0(hps_io_qspi_inst_IO2_0),
	.hps_io_qspi_inst_IO3_0(hps_io_qspi_inst_IO3_0),
	.hps_io_sdio_inst_CMD_0(hps_io_sdio_inst_CMD_0),
	.hps_io_sdio_inst_D0_0(hps_io_sdio_inst_D0_0),
	.hps_io_sdio_inst_D1_0(hps_io_sdio_inst_D1_0),
	.hps_io_sdio_inst_D2_0(hps_io_sdio_inst_D2_0),
	.hps_io_sdio_inst_D3_0(hps_io_sdio_inst_D3_0),
	.hps_io_usb1_inst_D0_0(hps_io_usb1_inst_D0_0),
	.hps_io_usb1_inst_D1_0(hps_io_usb1_inst_D1_0),
	.hps_io_usb1_inst_D2_0(hps_io_usb1_inst_D2_0),
	.hps_io_usb1_inst_D3_0(hps_io_usb1_inst_D3_0),
	.hps_io_usb1_inst_D4_0(hps_io_usb1_inst_D4_0),
	.hps_io_usb1_inst_D5_0(hps_io_usb1_inst_D5_0),
	.hps_io_usb1_inst_D6_0(hps_io_usb1_inst_D6_0),
	.hps_io_usb1_inst_D7_0(hps_io_usb1_inst_D7_0),
	.hps_io_i2c0_inst_SDA_0(hps_io_i2c0_inst_SDA_0),
	.hps_io_i2c0_inst_SCL_0(hps_io_i2c0_inst_SCL_0),
	.hps_io_i2c1_inst_SDA_0(hps_io_i2c1_inst_SDA_0),
	.hps_io_i2c1_inst_SCL_0(hps_io_i2c1_inst_SCL_0),
	.hps_io_gpio_inst_GPIO09_0(hps_io_gpio_inst_GPIO09_0),
	.hps_io_gpio_inst_GPIO35_0(hps_io_gpio_inst_GPIO35_0),
	.hps_io_gpio_inst_GPIO40_0(hps_io_gpio_inst_GPIO40_0),
	.hps_io_gpio_inst_GPIO41_0(hps_io_gpio_inst_GPIO41_0),
	.hps_io_gpio_inst_GPIO48_0(hps_io_gpio_inst_GPIO48_0),
	.hps_io_gpio_inst_GPIO53_0(hps_io_gpio_inst_GPIO53_0),
	.hps_io_gpio_inst_GPIO54_0(hps_io_gpio_inst_GPIO54_0),
	.hps_io_gpio_inst_GPIO61_0(hps_io_gpio_inst_GPIO61_0),
	.hps_io_hps_io_emac1_inst_RXD0(hps_io_hps_io_emac1_inst_RXD0),
	.hps_io_hps_io_emac1_inst_RXD1(hps_io_hps_io_emac1_inst_RXD1),
	.hps_io_hps_io_emac1_inst_RXD2(hps_io_hps_io_emac1_inst_RXD2),
	.hps_io_hps_io_emac1_inst_RXD3(hps_io_hps_io_emac1_inst_RXD3),
	.hps_io_hps_io_emac1_inst_RX_CLK(hps_io_hps_io_emac1_inst_RX_CLK),
	.hps_io_hps_io_emac1_inst_RX_CTL(hps_io_hps_io_emac1_inst_RX_CTL),
	.hps_io_hps_io_spim1_inst_MISO(hps_io_hps_io_spim1_inst_MISO),
	.hps_io_hps_io_uart0_inst_RX(hps_io_hps_io_uart0_inst_RX),
	.hps_io_hps_io_usb1_inst_CLK(hps_io_hps_io_usb1_inst_CLK),
	.hps_io_hps_io_usb1_inst_DIR(hps_io_hps_io_usb1_inst_DIR),
	.hps_io_hps_io_usb1_inst_NXT(hps_io_hps_io_usb1_inst_NXT),
	.memory_oct_rzqin(memory_oct_rzqin));

Computer_System_Computer_System_ARM_A9_HPS_fpga_interfaces fpga_interfaces(
	.h2f_rst_n({h2f_rst_n_0}),
	.h2f_lw_ARVALID({h2f_lw_ARVALID_0}),
	.h2f_lw_AWVALID({h2f_lw_AWVALID_0}),
	.h2f_lw_BREADY({h2f_lw_BREADY_0}),
	.h2f_lw_RREADY({h2f_lw_RREADY_0}),
	.h2f_lw_WLAST({h2f_lw_WLAST_0}),
	.h2f_lw_WVALID({h2f_lw_WVALID_0}),
	.h2f_lw_ARADDR({h2f_lw_ARADDR_unconnected_wire_20,h2f_lw_ARADDR_unconnected_wire_19,h2f_lw_ARADDR_unconnected_wire_18,h2f_lw_ARADDR_unconnected_wire_17,h2f_lw_ARADDR_unconnected_wire_16,h2f_lw_ARADDR_unconnected_wire_15,h2f_lw_ARADDR_unconnected_wire_14,
h2f_lw_ARADDR_unconnected_wire_13,h2f_lw_ARADDR_unconnected_wire_12,h2f_lw_ARADDR_unconnected_wire_11,h2f_lw_ARADDR_unconnected_wire_10,h2f_lw_ARADDR_unconnected_wire_9,h2f_lw_ARADDR_unconnected_wire_8,h2f_lw_ARADDR_unconnected_wire_7,
h2f_lw_ARADDR_unconnected_wire_6,h2f_lw_ARADDR_unconnected_wire_5,h2f_lw_ARADDR_4,h2f_lw_ARADDR_3,h2f_lw_ARADDR_2,h2f_lw_ARADDR_1,h2f_lw_ARADDR_0}),
	.h2f_lw_ARBURST({h2f_lw_ARBURST_1,h2f_lw_ARBURST_0}),
	.h2f_lw_ARID({h2f_lw_ARID_11,h2f_lw_ARID_10,h2f_lw_ARID_9,h2f_lw_ARID_8,h2f_lw_ARID_7,h2f_lw_ARID_6,h2f_lw_ARID_5,h2f_lw_ARID_4,h2f_lw_ARID_3,h2f_lw_ARID_2,h2f_lw_ARID_1,h2f_lw_ARID_0}),
	.h2f_lw_ARLEN({h2f_lw_ARLEN_3,h2f_lw_ARLEN_2,h2f_lw_ARLEN_1,h2f_lw_ARLEN_0}),
	.h2f_lw_ARSIZE({h2f_lw_ARSIZE_2,h2f_lw_ARSIZE_1,h2f_lw_ARSIZE_0}),
	.h2f_lw_AWADDR({h2f_lw_AWADDR_unconnected_wire_20,h2f_lw_AWADDR_unconnected_wire_19,h2f_lw_AWADDR_unconnected_wire_18,h2f_lw_AWADDR_unconnected_wire_17,h2f_lw_AWADDR_unconnected_wire_16,h2f_lw_AWADDR_unconnected_wire_15,h2f_lw_AWADDR_unconnected_wire_14,
h2f_lw_AWADDR_unconnected_wire_13,h2f_lw_AWADDR_unconnected_wire_12,h2f_lw_AWADDR_unconnected_wire_11,h2f_lw_AWADDR_unconnected_wire_10,h2f_lw_AWADDR_unconnected_wire_9,h2f_lw_AWADDR_unconnected_wire_8,h2f_lw_AWADDR_unconnected_wire_7,
h2f_lw_AWADDR_unconnected_wire_6,h2f_lw_AWADDR_unconnected_wire_5,h2f_lw_AWADDR_4,h2f_lw_AWADDR_3,h2f_lw_AWADDR_2,h2f_lw_AWADDR_1,h2f_lw_AWADDR_0}),
	.h2f_lw_AWBURST({h2f_lw_AWBURST_1,h2f_lw_AWBURST_0}),
	.h2f_lw_AWID({h2f_lw_AWID_11,h2f_lw_AWID_10,h2f_lw_AWID_9,h2f_lw_AWID_8,h2f_lw_AWID_7,h2f_lw_AWID_6,h2f_lw_AWID_5,h2f_lw_AWID_4,h2f_lw_AWID_3,h2f_lw_AWID_2,h2f_lw_AWID_1,h2f_lw_AWID_0}),
	.h2f_lw_AWLEN({h2f_lw_AWLEN_3,h2f_lw_AWLEN_2,h2f_lw_AWLEN_1,h2f_lw_AWLEN_0}),
	.h2f_lw_AWSIZE({h2f_lw_AWSIZE_2,h2f_lw_AWSIZE_1,h2f_lw_AWSIZE_0}),
	.h2f_lw_WDATA({h2f_lw_WDATA_31,h2f_lw_WDATA_30,h2f_lw_WDATA_29,h2f_lw_WDATA_28,h2f_lw_WDATA_27,h2f_lw_WDATA_26,h2f_lw_WDATA_25,h2f_lw_WDATA_24,h2f_lw_WDATA_23,h2f_lw_WDATA_22,h2f_lw_WDATA_21,h2f_lw_WDATA_20,h2f_lw_WDATA_19,h2f_lw_WDATA_18,h2f_lw_WDATA_17,h2f_lw_WDATA_16,h2f_lw_WDATA_15,
h2f_lw_WDATA_14,h2f_lw_WDATA_13,h2f_lw_WDATA_12,h2f_lw_WDATA_11,h2f_lw_WDATA_10,h2f_lw_WDATA_9,h2f_lw_WDATA_8,h2f_lw_WDATA_7,h2f_lw_WDATA_6,h2f_lw_WDATA_5,h2f_lw_WDATA_4,h2f_lw_WDATA_3,h2f_lw_WDATA_2,h2f_lw_WDATA_1,h2f_lw_WDATA_0}),
	.h2f_lw_WSTRB({h2f_lw_WSTRB_3,h2f_lw_WSTRB_2,h2f_lw_WSTRB_1,h2f_lw_WSTRB_0}),
	.h2f_ARVALID({h2f_ARVALID_0}),
	.h2f_AWVALID({h2f_AWVALID_0}),
	.h2f_BREADY({h2f_BREADY_0}),
	.h2f_RREADY({h2f_RREADY_0}),
	.h2f_WLAST({h2f_WLAST_0}),
	.h2f_WVALID({h2f_WVALID_0}),
	.h2f_ARADDR({h2f_ARADDR_unconnected_wire_29,h2f_ARADDR_unconnected_wire_28,h2f_ARADDR_unconnected_wire_27,h2f_ARADDR_unconnected_wire_26,h2f_ARADDR_unconnected_wire_25,h2f_ARADDR_unconnected_wire_24,h2f_ARADDR_unconnected_wire_23,h2f_ARADDR_unconnected_wire_22,
h2f_ARADDR_unconnected_wire_21,h2f_ARADDR_unconnected_wire_20,h2f_ARADDR_unconnected_wire_19,h2f_ARADDR_unconnected_wire_18,h2f_ARADDR_unconnected_wire_17,h2f_ARADDR_unconnected_wire_16,h2f_ARADDR_unconnected_wire_15,h2f_ARADDR_unconnected_wire_14,
h2f_ARADDR_unconnected_wire_13,h2f_ARADDR_unconnected_wire_12,h2f_ARADDR_unconnected_wire_11,h2f_ARADDR_unconnected_wire_10,h2f_ARADDR_9,h2f_ARADDR_8,h2f_ARADDR_7,h2f_ARADDR_6,h2f_ARADDR_5,h2f_ARADDR_4,h2f_ARADDR_3,h2f_ARADDR_2,h2f_ARADDR_1,h2f_ARADDR_0}),
	.h2f_ARBURST({h2f_ARBURST_1,h2f_ARBURST_0}),
	.h2f_ARID({h2f_ARID_11,h2f_ARID_10,h2f_ARID_9,h2f_ARID_8,h2f_ARID_7,h2f_ARID_6,h2f_ARID_5,h2f_ARID_4,h2f_ARID_3,h2f_ARID_2,h2f_ARID_1,h2f_ARID_0}),
	.h2f_ARLEN({h2f_ARLEN_3,h2f_ARLEN_2,h2f_ARLEN_1,h2f_ARLEN_0}),
	.h2f_ARSIZE({h2f_ARSIZE_2,h2f_ARSIZE_1,h2f_ARSIZE_0}),
	.h2f_AWADDR({h2f_AWADDR_unconnected_wire_29,h2f_AWADDR_unconnected_wire_28,h2f_AWADDR_27,h2f_AWADDR_26,h2f_AWADDR_25,h2f_AWADDR_24,h2f_AWADDR_23,h2f_AWADDR_22,h2f_AWADDR_21,h2f_AWADDR_20,h2f_AWADDR_19,h2f_AWADDR_18,h2f_AWADDR_17,h2f_AWADDR_16,h2f_AWADDR_15,h2f_AWADDR_14,h2f_AWADDR_13,
h2f_AWADDR_12,h2f_AWADDR_11,h2f_AWADDR_10,h2f_AWADDR_9,h2f_AWADDR_8,h2f_AWADDR_7,h2f_AWADDR_6,h2f_AWADDR_5,h2f_AWADDR_4,h2f_AWADDR_3,h2f_AWADDR_2,h2f_AWADDR_1,h2f_AWADDR_0}),
	.h2f_AWBURST({h2f_AWBURST_1,h2f_AWBURST_0}),
	.h2f_AWID({h2f_AWID_11,h2f_AWID_10,h2f_AWID_9,h2f_AWID_8,h2f_AWID_7,h2f_AWID_6,h2f_AWID_5,h2f_AWID_4,h2f_AWID_3,h2f_AWID_2,h2f_AWID_1,h2f_AWID_0}),
	.h2f_AWLEN({h2f_AWLEN_3,h2f_AWLEN_2,h2f_AWLEN_1,h2f_AWLEN_0}),
	.h2f_AWSIZE({h2f_AWSIZE_2,h2f_AWSIZE_1,h2f_AWSIZE_0}),
	.h2f_WDATA({h2f_WDATA_127,h2f_WDATA_126,h2f_WDATA_125,h2f_WDATA_124,h2f_WDATA_123,h2f_WDATA_122,h2f_WDATA_121,h2f_WDATA_120,h2f_WDATA_119,h2f_WDATA_118,h2f_WDATA_117,h2f_WDATA_116,h2f_WDATA_115,h2f_WDATA_114,h2f_WDATA_113,h2f_WDATA_112,h2f_WDATA_111,h2f_WDATA_110,h2f_WDATA_109,
h2f_WDATA_108,h2f_WDATA_107,h2f_WDATA_106,h2f_WDATA_105,h2f_WDATA_104,h2f_WDATA_103,h2f_WDATA_102,h2f_WDATA_101,h2f_WDATA_100,h2f_WDATA_99,h2f_WDATA_98,h2f_WDATA_97,h2f_WDATA_96,h2f_WDATA_95,h2f_WDATA_94,h2f_WDATA_93,h2f_WDATA_92,h2f_WDATA_91,h2f_WDATA_90,h2f_WDATA_89,
h2f_WDATA_88,h2f_WDATA_87,h2f_WDATA_86,h2f_WDATA_85,h2f_WDATA_84,h2f_WDATA_83,h2f_WDATA_82,h2f_WDATA_81,h2f_WDATA_80,h2f_WDATA_79,h2f_WDATA_78,h2f_WDATA_77,h2f_WDATA_76,h2f_WDATA_75,h2f_WDATA_74,h2f_WDATA_73,h2f_WDATA_72,h2f_WDATA_71,h2f_WDATA_70,h2f_WDATA_69,h2f_WDATA_68,
h2f_WDATA_67,h2f_WDATA_66,h2f_WDATA_65,h2f_WDATA_64,h2f_WDATA_63,h2f_WDATA_62,h2f_WDATA_61,h2f_WDATA_60,h2f_WDATA_59,h2f_WDATA_58,h2f_WDATA_57,h2f_WDATA_56,h2f_WDATA_55,h2f_WDATA_54,h2f_WDATA_53,h2f_WDATA_52,h2f_WDATA_51,h2f_WDATA_50,h2f_WDATA_49,h2f_WDATA_48,h2f_WDATA_47,
h2f_WDATA_46,h2f_WDATA_45,h2f_WDATA_44,h2f_WDATA_43,h2f_WDATA_42,h2f_WDATA_41,h2f_WDATA_40,h2f_WDATA_39,h2f_WDATA_38,h2f_WDATA_37,h2f_WDATA_36,h2f_WDATA_35,h2f_WDATA_34,h2f_WDATA_33,h2f_WDATA_32,h2f_WDATA_31,h2f_WDATA_30,h2f_WDATA_29,h2f_WDATA_28,h2f_WDATA_27,h2f_WDATA_26,
h2f_WDATA_25,h2f_WDATA_24,h2f_WDATA_23,h2f_WDATA_22,h2f_WDATA_21,h2f_WDATA_20,h2f_WDATA_19,h2f_WDATA_18,h2f_WDATA_17,h2f_WDATA_16,h2f_WDATA_15,h2f_WDATA_14,h2f_WDATA_13,h2f_WDATA_12,h2f_WDATA_11,h2f_WDATA_10,h2f_WDATA_9,h2f_WDATA_8,h2f_WDATA_7,h2f_WDATA_6,h2f_WDATA_5,
h2f_WDATA_4,h2f_WDATA_3,h2f_WDATA_2,h2f_WDATA_1,h2f_WDATA_0}),
	.h2f_WSTRB({h2f_WSTRB_15,h2f_WSTRB_14,h2f_WSTRB_13,h2f_WSTRB_12,h2f_WSTRB_11,h2f_WSTRB_10,h2f_WSTRB_9,h2f_WSTRB_8,h2f_WSTRB_7,h2f_WSTRB_6,h2f_WSTRB_5,h2f_WSTRB_4,h2f_WSTRB_3,h2f_WSTRB_2,h2f_WSTRB_1,h2f_WSTRB_0}),
	.h2f_lw_axi_clk({outclk_wire_0}),
	.f2h_axi_clk({outclk_wire_0}),
	.h2f_axi_clk({outclk_wire_0}),
	.h2f_lw_ARREADY({sink1_ready}),
	.h2f_lw_AWREADY({awready}),
	.h2f_lw_BVALID({src0_valid}),
	.h2f_lw_RLAST({source_endofpacket}),
	.h2f_lw_RVALID({src1_valid}),
	.h2f_lw_WREADY({wready}),
	.h2f_lw_BID({mem_99_0,mem_98_0,mem_97_0,mem_96_0,mem_95_0,mem_94_0,mem_93_0,mem_92_0,mem_91_0,mem_90_0,mem_89_0,mem_88_0}),
	.h2f_lw_RID({mem_99_0,mem_98_0,mem_97_0,mem_96_0,mem_95_0,mem_94_0,mem_93_0,mem_92_0,mem_91_0,mem_90_0,mem_89_0,mem_88_0}),
	.h2f_lw_RDATA({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,out_data_7,out_data_6,out_data_5,out_data_4,out_data_3,out_data_2,out_data_1,out_data_0}),
	.h2f_ARREADY({sink1_ready1}),
	.h2f_AWREADY({awready1}),
	.h2f_BVALID({WideOr1}),
	.h2f_RLAST({src_payload_0}),
	.h2f_RVALID({WideOr11}),
	.h2f_WREADY({wready1}),
	.h2f_BID({src_data_220,src_data_219,src_data_218,src_data_217,src_data_216,src_data_215,src_data_214,src_data_213,src_data_212,src_data_211,src_data_210,src_data_209}),
	.h2f_RDATA({src_data_127,src_data_126,src_payload39,src_data_124,src_data_123,src_data_122,src_data_121,src_payload38,src_data_119,src_payload37,src_data_117,src_payload36,src_data_115,src_data_114,src_payload35,src_data_112,src_data_111,src_data_110,src_payload34,src_data_108,
src_data_107,src_data_106,src_data_105,src_payload33,src_data_103,src_payload32,src_data_101,src_payload31,src_data_99,src_data_98,src_payload30,src_data_96,src_data_95,src_data_94,src_payload29,src_data_92,src_data_91,src_data_90,src_data_89,src_payload28,src_data_87,
src_payload27,src_data_85,src_payload26,src_data_83,src_data_82,src_payload25,src_data_80,src_data_79,src_data_78,src_payload24,src_data_76,src_data_75,src_data_74,src_data_73,src_payload23,src_data_71,src_payload22,src_data_69,src_payload21,src_data_67,src_data_66,
src_payload20,src_data_64,src_data_63,src_data_62,src_payload19,src_data_60,src_data_59,src_data_58,src_data_57,src_payload18,src_data_55,src_payload17,src_data_53,src_payload16,src_data_51,src_data_50,src_payload15,src_data_48,src_data_47,src_data_46,src_payload14,src_data_44,
src_data_43,src_data_42,src_data_41,src_payload13,src_data_39,src_payload12,src_data_37,src_payload11,src_data_35,src_data_34,src_payload10,src_data_32,src_data_31,src_data_30,src_payload9,src_data_28,src_data_27,src_data_26,src_data_25,src_payload8,src_data_23,src_payload7,
src_data_21,src_payload6,src_data_19,src_data_18,src_payload5,src_data_16,src_data_15,src_data_14,src_payload4,src_data_12,src_data_11,src_data_10,src_data_9,src_payload3,src_data_7,src_payload2,src_data_5,src_payload1,src_data_3,src_data_2,src_payload,src_data_0}),
	.h2f_RID({src_data_2201,src_data_2191,src_data_2181,src_data_2171,src_data_2161,src_data_2151,src_data_2141,src_data_2131,src_data_2121,src_data_2111,src_data_2101,src_data_2091}));

endmodule

module Computer_System_Computer_System_ARM_A9_HPS_fpga_interfaces (
	h2f_rst_n,
	h2f_lw_ARVALID,
	h2f_lw_AWVALID,
	h2f_lw_BREADY,
	h2f_lw_RREADY,
	h2f_lw_WLAST,
	h2f_lw_WVALID,
	h2f_lw_ARADDR,
	h2f_lw_ARBURST,
	h2f_lw_ARID,
	h2f_lw_ARLEN,
	h2f_lw_ARSIZE,
	h2f_lw_AWADDR,
	h2f_lw_AWBURST,
	h2f_lw_AWID,
	h2f_lw_AWLEN,
	h2f_lw_AWSIZE,
	h2f_lw_WDATA,
	h2f_lw_WSTRB,
	h2f_ARVALID,
	h2f_AWVALID,
	h2f_BREADY,
	h2f_RREADY,
	h2f_WLAST,
	h2f_WVALID,
	h2f_ARADDR,
	h2f_ARBURST,
	h2f_ARID,
	h2f_ARLEN,
	h2f_ARSIZE,
	h2f_AWADDR,
	h2f_AWBURST,
	h2f_AWID,
	h2f_AWLEN,
	h2f_AWSIZE,
	h2f_WDATA,
	h2f_WSTRB,
	h2f_lw_axi_clk,
	f2h_axi_clk,
	h2f_axi_clk,
	h2f_lw_ARREADY,
	h2f_lw_AWREADY,
	h2f_lw_BVALID,
	h2f_lw_RLAST,
	h2f_lw_RVALID,
	h2f_lw_WREADY,
	h2f_lw_BID,
	h2f_lw_RID,
	h2f_lw_RDATA,
	h2f_ARREADY,
	h2f_AWREADY,
	h2f_BVALID,
	h2f_RLAST,
	h2f_RVALID,
	h2f_WREADY,
	h2f_BID,
	h2f_RDATA,
	h2f_RID)/* synthesis synthesis_greybox=0 */;
output 	[0:0] h2f_rst_n;
output 	[0:0] h2f_lw_ARVALID;
output 	[0:0] h2f_lw_AWVALID;
output 	[0:0] h2f_lw_BREADY;
output 	[0:0] h2f_lw_RREADY;
output 	[0:0] h2f_lw_WLAST;
output 	[0:0] h2f_lw_WVALID;
output 	[20:0] h2f_lw_ARADDR;
output 	[1:0] h2f_lw_ARBURST;
output 	[11:0] h2f_lw_ARID;
output 	[3:0] h2f_lw_ARLEN;
output 	[2:0] h2f_lw_ARSIZE;
output 	[20:0] h2f_lw_AWADDR;
output 	[1:0] h2f_lw_AWBURST;
output 	[11:0] h2f_lw_AWID;
output 	[3:0] h2f_lw_AWLEN;
output 	[2:0] h2f_lw_AWSIZE;
output 	[31:0] h2f_lw_WDATA;
output 	[3:0] h2f_lw_WSTRB;
output 	[0:0] h2f_ARVALID;
output 	[0:0] h2f_AWVALID;
output 	[0:0] h2f_BREADY;
output 	[0:0] h2f_RREADY;
output 	[0:0] h2f_WLAST;
output 	[0:0] h2f_WVALID;
output 	[29:0] h2f_ARADDR;
output 	[1:0] h2f_ARBURST;
output 	[11:0] h2f_ARID;
output 	[3:0] h2f_ARLEN;
output 	[2:0] h2f_ARSIZE;
output 	[29:0] h2f_AWADDR;
output 	[1:0] h2f_AWBURST;
output 	[11:0] h2f_AWID;
output 	[3:0] h2f_AWLEN;
output 	[2:0] h2f_AWSIZE;
output 	[127:0] h2f_WDATA;
output 	[15:0] h2f_WSTRB;
input 	[0:0] h2f_lw_axi_clk;
input 	[0:0] f2h_axi_clk;
input 	[0:0] h2f_axi_clk;
input 	[0:0] h2f_lw_ARREADY;
input 	[0:0] h2f_lw_AWREADY;
input 	[0:0] h2f_lw_BVALID;
input 	[0:0] h2f_lw_RLAST;
input 	[0:0] h2f_lw_RVALID;
input 	[0:0] h2f_lw_WREADY;
input 	[11:0] h2f_lw_BID;
input 	[11:0] h2f_lw_RID;
input 	[31:0] h2f_lw_RDATA;
input 	[0:0] h2f_ARREADY;
input 	[0:0] h2f_AWREADY;
input 	[0:0] h2f_BVALID;
input 	[0:0] h2f_RLAST;
input 	[0:0] h2f_RVALID;
input 	[0:0] h2f_WREADY;
input 	[11:0] h2f_BID;
input 	[127:0] h2f_RDATA;
input 	[11:0] h2f_RID;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \debug_apb~O_P_ADDR_31 ;
wire \tpiu~trace_data ;
wire \tpiu~O_TRACE_DATA1 ;
wire \tpiu~O_TRACE_DATA2 ;
wire \tpiu~O_TRACE_DATA3 ;
wire \tpiu~O_TRACE_DATA4 ;
wire \tpiu~O_TRACE_DATA5 ;
wire \tpiu~O_TRACE_DATA6 ;
wire \tpiu~O_TRACE_DATA7 ;
wire \tpiu~O_TRACE_DATA8 ;
wire \tpiu~O_TRACE_DATA9 ;
wire \tpiu~O_TRACE_DATA10 ;
wire \tpiu~O_TRACE_DATA11 ;
wire \tpiu~O_TRACE_DATA12 ;
wire \tpiu~O_TRACE_DATA13 ;
wire \tpiu~O_TRACE_DATA14 ;
wire \tpiu~O_TRACE_DATA15 ;
wire \tpiu~O_TRACE_DATA16 ;
wire \tpiu~O_TRACE_DATA17 ;
wire \tpiu~O_TRACE_DATA18 ;
wire \tpiu~O_TRACE_DATA19 ;
wire \tpiu~O_TRACE_DATA20 ;
wire \tpiu~O_TRACE_DATA21 ;
wire \tpiu~O_TRACE_DATA22 ;
wire \tpiu~O_TRACE_DATA23 ;
wire \tpiu~O_TRACE_DATA24 ;
wire \tpiu~O_TRACE_DATA25 ;
wire \tpiu~O_TRACE_DATA26 ;
wire \tpiu~O_TRACE_DATA27 ;
wire \tpiu~O_TRACE_DATA28 ;
wire \tpiu~O_TRACE_DATA29 ;
wire \tpiu~O_TRACE_DATA30 ;
wire \tpiu~O_TRACE_DATA31 ;
wire \boot_from_fpga~fake_dout ;
wire \f2h_ARREADY[0] ;
wire \f2sdram~O_BONDING_OUT_10 ;
wire \f2sdram~O_BONDING_OUT_11 ;
wire \f2sdram~O_BONDING_OUT_12 ;
wire \f2sdram~O_BONDING_OUT_13 ;
wire \interrupts~fake_dout ;
wire \clocks_resets~h2f_cold_rst_n ;
wire \h2f_lw_ARADDR[5] ;
wire \h2f_lw_ARADDR[6] ;
wire \h2f_lw_ARADDR[7] ;
wire \h2f_lw_ARADDR[8] ;
wire \h2f_lw_ARADDR[9] ;
wire \h2f_lw_ARADDR[10] ;
wire \h2f_lw_ARADDR[11] ;
wire \h2f_lw_ARADDR[12] ;
wire \h2f_lw_ARADDR[13] ;
wire \h2f_lw_ARADDR[14] ;
wire \h2f_lw_ARADDR[15] ;
wire \h2f_lw_ARADDR[16] ;
wire \h2f_lw_ARADDR[17] ;
wire \h2f_lw_ARADDR[18] ;
wire \h2f_lw_ARADDR[19] ;
wire \h2f_lw_ARADDR[20] ;
wire \h2f_ARADDR[10] ;
wire \h2f_ARADDR[11] ;
wire \h2f_ARADDR[12] ;
wire \h2f_ARADDR[13] ;
wire \h2f_ARADDR[14] ;
wire \h2f_ARADDR[15] ;
wire \h2f_ARADDR[16] ;
wire \h2f_ARADDR[17] ;
wire \h2f_ARADDR[18] ;
wire \h2f_ARADDR[19] ;
wire \h2f_ARADDR[20] ;
wire \h2f_ARADDR[21] ;
wire \h2f_ARADDR[22] ;
wire \h2f_ARADDR[23] ;
wire \h2f_ARADDR[24] ;
wire \h2f_ARADDR[25] ;
wire \h2f_ARADDR[26] ;
wire \h2f_ARADDR[27] ;
wire \h2f_ARADDR[28] ;
wire \h2f_ARADDR[29] ;

wire [31:0] tpiu_TRACE_DATA_bus;
wire [3:0] f2sdram_BONDING_OUT_1_bus;
wire [20:0] hps2fpga_light_weight_ARADDR_bus;
wire [1:0] hps2fpga_light_weight_ARBURST_bus;
wire [11:0] hps2fpga_light_weight_ARID_bus;
wire [3:0] hps2fpga_light_weight_ARLEN_bus;
wire [2:0] hps2fpga_light_weight_ARSIZE_bus;
wire [20:0] hps2fpga_light_weight_AWADDR_bus;
wire [1:0] hps2fpga_light_weight_AWBURST_bus;
wire [11:0] hps2fpga_light_weight_AWID_bus;
wire [3:0] hps2fpga_light_weight_AWLEN_bus;
wire [2:0] hps2fpga_light_weight_AWSIZE_bus;
wire [31:0] hps2fpga_light_weight_WDATA_bus;
wire [3:0] hps2fpga_light_weight_WSTRB_bus;
wire [29:0] hps2fpga_ARADDR_bus;
wire [1:0] hps2fpga_ARBURST_bus;
wire [11:0] hps2fpga_ARID_bus;
wire [3:0] hps2fpga_ARLEN_bus;
wire [2:0] hps2fpga_ARSIZE_bus;
wire [29:0] hps2fpga_AWADDR_bus;
wire [1:0] hps2fpga_AWBURST_bus;
wire [11:0] hps2fpga_AWID_bus;
wire [3:0] hps2fpga_AWLEN_bus;
wire [2:0] hps2fpga_AWSIZE_bus;
wire [127:0] hps2fpga_WDATA_bus;
wire [15:0] hps2fpga_WSTRB_bus;

assign \tpiu~trace_data  = tpiu_TRACE_DATA_bus[0];
assign \tpiu~O_TRACE_DATA1  = tpiu_TRACE_DATA_bus[1];
assign \tpiu~O_TRACE_DATA2  = tpiu_TRACE_DATA_bus[2];
assign \tpiu~O_TRACE_DATA3  = tpiu_TRACE_DATA_bus[3];
assign \tpiu~O_TRACE_DATA4  = tpiu_TRACE_DATA_bus[4];
assign \tpiu~O_TRACE_DATA5  = tpiu_TRACE_DATA_bus[5];
assign \tpiu~O_TRACE_DATA6  = tpiu_TRACE_DATA_bus[6];
assign \tpiu~O_TRACE_DATA7  = tpiu_TRACE_DATA_bus[7];
assign \tpiu~O_TRACE_DATA8  = tpiu_TRACE_DATA_bus[8];
assign \tpiu~O_TRACE_DATA9  = tpiu_TRACE_DATA_bus[9];
assign \tpiu~O_TRACE_DATA10  = tpiu_TRACE_DATA_bus[10];
assign \tpiu~O_TRACE_DATA11  = tpiu_TRACE_DATA_bus[11];
assign \tpiu~O_TRACE_DATA12  = tpiu_TRACE_DATA_bus[12];
assign \tpiu~O_TRACE_DATA13  = tpiu_TRACE_DATA_bus[13];
assign \tpiu~O_TRACE_DATA14  = tpiu_TRACE_DATA_bus[14];
assign \tpiu~O_TRACE_DATA15  = tpiu_TRACE_DATA_bus[15];
assign \tpiu~O_TRACE_DATA16  = tpiu_TRACE_DATA_bus[16];
assign \tpiu~O_TRACE_DATA17  = tpiu_TRACE_DATA_bus[17];
assign \tpiu~O_TRACE_DATA18  = tpiu_TRACE_DATA_bus[18];
assign \tpiu~O_TRACE_DATA19  = tpiu_TRACE_DATA_bus[19];
assign \tpiu~O_TRACE_DATA20  = tpiu_TRACE_DATA_bus[20];
assign \tpiu~O_TRACE_DATA21  = tpiu_TRACE_DATA_bus[21];
assign \tpiu~O_TRACE_DATA22  = tpiu_TRACE_DATA_bus[22];
assign \tpiu~O_TRACE_DATA23  = tpiu_TRACE_DATA_bus[23];
assign \tpiu~O_TRACE_DATA24  = tpiu_TRACE_DATA_bus[24];
assign \tpiu~O_TRACE_DATA25  = tpiu_TRACE_DATA_bus[25];
assign \tpiu~O_TRACE_DATA26  = tpiu_TRACE_DATA_bus[26];
assign \tpiu~O_TRACE_DATA27  = tpiu_TRACE_DATA_bus[27];
assign \tpiu~O_TRACE_DATA28  = tpiu_TRACE_DATA_bus[28];
assign \tpiu~O_TRACE_DATA29  = tpiu_TRACE_DATA_bus[29];
assign \tpiu~O_TRACE_DATA30  = tpiu_TRACE_DATA_bus[30];
assign \tpiu~O_TRACE_DATA31  = tpiu_TRACE_DATA_bus[31];

assign \f2sdram~O_BONDING_OUT_10  = f2sdram_BONDING_OUT_1_bus[0];
assign \f2sdram~O_BONDING_OUT_11  = f2sdram_BONDING_OUT_1_bus[1];
assign \f2sdram~O_BONDING_OUT_12  = f2sdram_BONDING_OUT_1_bus[2];
assign \f2sdram~O_BONDING_OUT_13  = f2sdram_BONDING_OUT_1_bus[3];

assign h2f_lw_ARADDR[0] = hps2fpga_light_weight_ARADDR_bus[0];
assign h2f_lw_ARADDR[1] = hps2fpga_light_weight_ARADDR_bus[1];
assign h2f_lw_ARADDR[2] = hps2fpga_light_weight_ARADDR_bus[2];
assign h2f_lw_ARADDR[3] = hps2fpga_light_weight_ARADDR_bus[3];
assign h2f_lw_ARADDR[4] = hps2fpga_light_weight_ARADDR_bus[4];
assign \h2f_lw_ARADDR[5]  = hps2fpga_light_weight_ARADDR_bus[5];
assign \h2f_lw_ARADDR[6]  = hps2fpga_light_weight_ARADDR_bus[6];
assign \h2f_lw_ARADDR[7]  = hps2fpga_light_weight_ARADDR_bus[7];
assign \h2f_lw_ARADDR[8]  = hps2fpga_light_weight_ARADDR_bus[8];
assign \h2f_lw_ARADDR[9]  = hps2fpga_light_weight_ARADDR_bus[9];
assign \h2f_lw_ARADDR[10]  = hps2fpga_light_weight_ARADDR_bus[10];
assign \h2f_lw_ARADDR[11]  = hps2fpga_light_weight_ARADDR_bus[11];
assign \h2f_lw_ARADDR[12]  = hps2fpga_light_weight_ARADDR_bus[12];
assign \h2f_lw_ARADDR[13]  = hps2fpga_light_weight_ARADDR_bus[13];
assign \h2f_lw_ARADDR[14]  = hps2fpga_light_weight_ARADDR_bus[14];
assign \h2f_lw_ARADDR[15]  = hps2fpga_light_weight_ARADDR_bus[15];
assign \h2f_lw_ARADDR[16]  = hps2fpga_light_weight_ARADDR_bus[16];
assign \h2f_lw_ARADDR[17]  = hps2fpga_light_weight_ARADDR_bus[17];
assign \h2f_lw_ARADDR[18]  = hps2fpga_light_weight_ARADDR_bus[18];
assign \h2f_lw_ARADDR[19]  = hps2fpga_light_weight_ARADDR_bus[19];
assign \h2f_lw_ARADDR[20]  = hps2fpga_light_weight_ARADDR_bus[20];

assign h2f_lw_ARBURST[0] = hps2fpga_light_weight_ARBURST_bus[0];
assign h2f_lw_ARBURST[1] = hps2fpga_light_weight_ARBURST_bus[1];

assign h2f_lw_ARID[0] = hps2fpga_light_weight_ARID_bus[0];
assign h2f_lw_ARID[1] = hps2fpga_light_weight_ARID_bus[1];
assign h2f_lw_ARID[2] = hps2fpga_light_weight_ARID_bus[2];
assign h2f_lw_ARID[3] = hps2fpga_light_weight_ARID_bus[3];
assign h2f_lw_ARID[4] = hps2fpga_light_weight_ARID_bus[4];
assign h2f_lw_ARID[5] = hps2fpga_light_weight_ARID_bus[5];
assign h2f_lw_ARID[6] = hps2fpga_light_weight_ARID_bus[6];
assign h2f_lw_ARID[7] = hps2fpga_light_weight_ARID_bus[7];
assign h2f_lw_ARID[8] = hps2fpga_light_weight_ARID_bus[8];
assign h2f_lw_ARID[9] = hps2fpga_light_weight_ARID_bus[9];
assign h2f_lw_ARID[10] = hps2fpga_light_weight_ARID_bus[10];
assign h2f_lw_ARID[11] = hps2fpga_light_weight_ARID_bus[11];

assign h2f_lw_ARLEN[0] = hps2fpga_light_weight_ARLEN_bus[0];
assign h2f_lw_ARLEN[1] = hps2fpga_light_weight_ARLEN_bus[1];
assign h2f_lw_ARLEN[2] = hps2fpga_light_weight_ARLEN_bus[2];
assign h2f_lw_ARLEN[3] = hps2fpga_light_weight_ARLEN_bus[3];

assign h2f_lw_ARSIZE[0] = hps2fpga_light_weight_ARSIZE_bus[0];
assign h2f_lw_ARSIZE[1] = hps2fpga_light_weight_ARSIZE_bus[1];
assign h2f_lw_ARSIZE[2] = hps2fpga_light_weight_ARSIZE_bus[2];

assign h2f_lw_AWADDR[0] = hps2fpga_light_weight_AWADDR_bus[0];
assign h2f_lw_AWADDR[1] = hps2fpga_light_weight_AWADDR_bus[1];
assign h2f_lw_AWADDR[2] = hps2fpga_light_weight_AWADDR_bus[2];
assign h2f_lw_AWADDR[3] = hps2fpga_light_weight_AWADDR_bus[3];
assign h2f_lw_AWADDR[4] = hps2fpga_light_weight_AWADDR_bus[4];

assign h2f_lw_AWBURST[0] = hps2fpga_light_weight_AWBURST_bus[0];
assign h2f_lw_AWBURST[1] = hps2fpga_light_weight_AWBURST_bus[1];

assign h2f_lw_AWID[0] = hps2fpga_light_weight_AWID_bus[0];
assign h2f_lw_AWID[1] = hps2fpga_light_weight_AWID_bus[1];
assign h2f_lw_AWID[2] = hps2fpga_light_weight_AWID_bus[2];
assign h2f_lw_AWID[3] = hps2fpga_light_weight_AWID_bus[3];
assign h2f_lw_AWID[4] = hps2fpga_light_weight_AWID_bus[4];
assign h2f_lw_AWID[5] = hps2fpga_light_weight_AWID_bus[5];
assign h2f_lw_AWID[6] = hps2fpga_light_weight_AWID_bus[6];
assign h2f_lw_AWID[7] = hps2fpga_light_weight_AWID_bus[7];
assign h2f_lw_AWID[8] = hps2fpga_light_weight_AWID_bus[8];
assign h2f_lw_AWID[9] = hps2fpga_light_weight_AWID_bus[9];
assign h2f_lw_AWID[10] = hps2fpga_light_weight_AWID_bus[10];
assign h2f_lw_AWID[11] = hps2fpga_light_weight_AWID_bus[11];

assign h2f_lw_AWLEN[0] = hps2fpga_light_weight_AWLEN_bus[0];
assign h2f_lw_AWLEN[1] = hps2fpga_light_weight_AWLEN_bus[1];
assign h2f_lw_AWLEN[2] = hps2fpga_light_weight_AWLEN_bus[2];
assign h2f_lw_AWLEN[3] = hps2fpga_light_weight_AWLEN_bus[3];

assign h2f_lw_AWSIZE[0] = hps2fpga_light_weight_AWSIZE_bus[0];
assign h2f_lw_AWSIZE[1] = hps2fpga_light_weight_AWSIZE_bus[1];
assign h2f_lw_AWSIZE[2] = hps2fpga_light_weight_AWSIZE_bus[2];

assign h2f_lw_WDATA[0] = hps2fpga_light_weight_WDATA_bus[0];
assign h2f_lw_WDATA[1] = hps2fpga_light_weight_WDATA_bus[1];
assign h2f_lw_WDATA[2] = hps2fpga_light_weight_WDATA_bus[2];
assign h2f_lw_WDATA[3] = hps2fpga_light_weight_WDATA_bus[3];
assign h2f_lw_WDATA[4] = hps2fpga_light_weight_WDATA_bus[4];
assign h2f_lw_WDATA[5] = hps2fpga_light_weight_WDATA_bus[5];
assign h2f_lw_WDATA[6] = hps2fpga_light_weight_WDATA_bus[6];
assign h2f_lw_WDATA[7] = hps2fpga_light_weight_WDATA_bus[7];
assign h2f_lw_WDATA[8] = hps2fpga_light_weight_WDATA_bus[8];
assign h2f_lw_WDATA[9] = hps2fpga_light_weight_WDATA_bus[9];
assign h2f_lw_WDATA[10] = hps2fpga_light_weight_WDATA_bus[10];
assign h2f_lw_WDATA[11] = hps2fpga_light_weight_WDATA_bus[11];
assign h2f_lw_WDATA[12] = hps2fpga_light_weight_WDATA_bus[12];
assign h2f_lw_WDATA[13] = hps2fpga_light_weight_WDATA_bus[13];
assign h2f_lw_WDATA[14] = hps2fpga_light_weight_WDATA_bus[14];
assign h2f_lw_WDATA[15] = hps2fpga_light_weight_WDATA_bus[15];
assign h2f_lw_WDATA[16] = hps2fpga_light_weight_WDATA_bus[16];
assign h2f_lw_WDATA[17] = hps2fpga_light_weight_WDATA_bus[17];
assign h2f_lw_WDATA[18] = hps2fpga_light_weight_WDATA_bus[18];
assign h2f_lw_WDATA[19] = hps2fpga_light_weight_WDATA_bus[19];
assign h2f_lw_WDATA[20] = hps2fpga_light_weight_WDATA_bus[20];
assign h2f_lw_WDATA[21] = hps2fpga_light_weight_WDATA_bus[21];
assign h2f_lw_WDATA[22] = hps2fpga_light_weight_WDATA_bus[22];
assign h2f_lw_WDATA[23] = hps2fpga_light_weight_WDATA_bus[23];
assign h2f_lw_WDATA[24] = hps2fpga_light_weight_WDATA_bus[24];
assign h2f_lw_WDATA[25] = hps2fpga_light_weight_WDATA_bus[25];
assign h2f_lw_WDATA[26] = hps2fpga_light_weight_WDATA_bus[26];
assign h2f_lw_WDATA[27] = hps2fpga_light_weight_WDATA_bus[27];
assign h2f_lw_WDATA[28] = hps2fpga_light_weight_WDATA_bus[28];
assign h2f_lw_WDATA[29] = hps2fpga_light_weight_WDATA_bus[29];
assign h2f_lw_WDATA[30] = hps2fpga_light_weight_WDATA_bus[30];
assign h2f_lw_WDATA[31] = hps2fpga_light_weight_WDATA_bus[31];

assign h2f_lw_WSTRB[0] = hps2fpga_light_weight_WSTRB_bus[0];
assign h2f_lw_WSTRB[1] = hps2fpga_light_weight_WSTRB_bus[1];
assign h2f_lw_WSTRB[2] = hps2fpga_light_weight_WSTRB_bus[2];
assign h2f_lw_WSTRB[3] = hps2fpga_light_weight_WSTRB_bus[3];

assign h2f_ARADDR[0] = hps2fpga_ARADDR_bus[0];
assign h2f_ARADDR[1] = hps2fpga_ARADDR_bus[1];
assign h2f_ARADDR[2] = hps2fpga_ARADDR_bus[2];
assign h2f_ARADDR[3] = hps2fpga_ARADDR_bus[3];
assign h2f_ARADDR[4] = hps2fpga_ARADDR_bus[4];
assign h2f_ARADDR[5] = hps2fpga_ARADDR_bus[5];
assign h2f_ARADDR[6] = hps2fpga_ARADDR_bus[6];
assign h2f_ARADDR[7] = hps2fpga_ARADDR_bus[7];
assign h2f_ARADDR[8] = hps2fpga_ARADDR_bus[8];
assign h2f_ARADDR[9] = hps2fpga_ARADDR_bus[9];
assign \h2f_ARADDR[10]  = hps2fpga_ARADDR_bus[10];
assign \h2f_ARADDR[11]  = hps2fpga_ARADDR_bus[11];
assign \h2f_ARADDR[12]  = hps2fpga_ARADDR_bus[12];
assign \h2f_ARADDR[13]  = hps2fpga_ARADDR_bus[13];
assign \h2f_ARADDR[14]  = hps2fpga_ARADDR_bus[14];
assign \h2f_ARADDR[15]  = hps2fpga_ARADDR_bus[15];
assign \h2f_ARADDR[16]  = hps2fpga_ARADDR_bus[16];
assign \h2f_ARADDR[17]  = hps2fpga_ARADDR_bus[17];
assign \h2f_ARADDR[18]  = hps2fpga_ARADDR_bus[18];
assign \h2f_ARADDR[19]  = hps2fpga_ARADDR_bus[19];
assign \h2f_ARADDR[20]  = hps2fpga_ARADDR_bus[20];
assign \h2f_ARADDR[21]  = hps2fpga_ARADDR_bus[21];
assign \h2f_ARADDR[22]  = hps2fpga_ARADDR_bus[22];
assign \h2f_ARADDR[23]  = hps2fpga_ARADDR_bus[23];
assign \h2f_ARADDR[24]  = hps2fpga_ARADDR_bus[24];
assign \h2f_ARADDR[25]  = hps2fpga_ARADDR_bus[25];
assign \h2f_ARADDR[26]  = hps2fpga_ARADDR_bus[26];
assign \h2f_ARADDR[27]  = hps2fpga_ARADDR_bus[27];
assign \h2f_ARADDR[28]  = hps2fpga_ARADDR_bus[28];
assign \h2f_ARADDR[29]  = hps2fpga_ARADDR_bus[29];

assign h2f_ARBURST[0] = hps2fpga_ARBURST_bus[0];
assign h2f_ARBURST[1] = hps2fpga_ARBURST_bus[1];

assign h2f_ARID[0] = hps2fpga_ARID_bus[0];
assign h2f_ARID[1] = hps2fpga_ARID_bus[1];
assign h2f_ARID[2] = hps2fpga_ARID_bus[2];
assign h2f_ARID[3] = hps2fpga_ARID_bus[3];
assign h2f_ARID[4] = hps2fpga_ARID_bus[4];
assign h2f_ARID[5] = hps2fpga_ARID_bus[5];
assign h2f_ARID[6] = hps2fpga_ARID_bus[6];
assign h2f_ARID[7] = hps2fpga_ARID_bus[7];
assign h2f_ARID[8] = hps2fpga_ARID_bus[8];
assign h2f_ARID[9] = hps2fpga_ARID_bus[9];
assign h2f_ARID[10] = hps2fpga_ARID_bus[10];
assign h2f_ARID[11] = hps2fpga_ARID_bus[11];

assign h2f_ARLEN[0] = hps2fpga_ARLEN_bus[0];
assign h2f_ARLEN[1] = hps2fpga_ARLEN_bus[1];
assign h2f_ARLEN[2] = hps2fpga_ARLEN_bus[2];
assign h2f_ARLEN[3] = hps2fpga_ARLEN_bus[3];

assign h2f_ARSIZE[0] = hps2fpga_ARSIZE_bus[0];
assign h2f_ARSIZE[1] = hps2fpga_ARSIZE_bus[1];
assign h2f_ARSIZE[2] = hps2fpga_ARSIZE_bus[2];

assign h2f_AWADDR[0] = hps2fpga_AWADDR_bus[0];
assign h2f_AWADDR[1] = hps2fpga_AWADDR_bus[1];
assign h2f_AWADDR[2] = hps2fpga_AWADDR_bus[2];
assign h2f_AWADDR[3] = hps2fpga_AWADDR_bus[3];
assign h2f_AWADDR[4] = hps2fpga_AWADDR_bus[4];
assign h2f_AWADDR[5] = hps2fpga_AWADDR_bus[5];
assign h2f_AWADDR[6] = hps2fpga_AWADDR_bus[6];
assign h2f_AWADDR[7] = hps2fpga_AWADDR_bus[7];
assign h2f_AWADDR[8] = hps2fpga_AWADDR_bus[8];
assign h2f_AWADDR[9] = hps2fpga_AWADDR_bus[9];
assign h2f_AWADDR[10] = hps2fpga_AWADDR_bus[10];
assign h2f_AWADDR[11] = hps2fpga_AWADDR_bus[11];
assign h2f_AWADDR[12] = hps2fpga_AWADDR_bus[12];
assign h2f_AWADDR[13] = hps2fpga_AWADDR_bus[13];
assign h2f_AWADDR[14] = hps2fpga_AWADDR_bus[14];
assign h2f_AWADDR[15] = hps2fpga_AWADDR_bus[15];
assign h2f_AWADDR[16] = hps2fpga_AWADDR_bus[16];
assign h2f_AWADDR[17] = hps2fpga_AWADDR_bus[17];
assign h2f_AWADDR[18] = hps2fpga_AWADDR_bus[18];
assign h2f_AWADDR[19] = hps2fpga_AWADDR_bus[19];
assign h2f_AWADDR[20] = hps2fpga_AWADDR_bus[20];
assign h2f_AWADDR[21] = hps2fpga_AWADDR_bus[21];
assign h2f_AWADDR[22] = hps2fpga_AWADDR_bus[22];
assign h2f_AWADDR[23] = hps2fpga_AWADDR_bus[23];
assign h2f_AWADDR[24] = hps2fpga_AWADDR_bus[24];
assign h2f_AWADDR[25] = hps2fpga_AWADDR_bus[25];
assign h2f_AWADDR[26] = hps2fpga_AWADDR_bus[26];
assign h2f_AWADDR[27] = hps2fpga_AWADDR_bus[27];

assign h2f_AWBURST[0] = hps2fpga_AWBURST_bus[0];
assign h2f_AWBURST[1] = hps2fpga_AWBURST_bus[1];

assign h2f_AWID[0] = hps2fpga_AWID_bus[0];
assign h2f_AWID[1] = hps2fpga_AWID_bus[1];
assign h2f_AWID[2] = hps2fpga_AWID_bus[2];
assign h2f_AWID[3] = hps2fpga_AWID_bus[3];
assign h2f_AWID[4] = hps2fpga_AWID_bus[4];
assign h2f_AWID[5] = hps2fpga_AWID_bus[5];
assign h2f_AWID[6] = hps2fpga_AWID_bus[6];
assign h2f_AWID[7] = hps2fpga_AWID_bus[7];
assign h2f_AWID[8] = hps2fpga_AWID_bus[8];
assign h2f_AWID[9] = hps2fpga_AWID_bus[9];
assign h2f_AWID[10] = hps2fpga_AWID_bus[10];
assign h2f_AWID[11] = hps2fpga_AWID_bus[11];

assign h2f_AWLEN[0] = hps2fpga_AWLEN_bus[0];
assign h2f_AWLEN[1] = hps2fpga_AWLEN_bus[1];
assign h2f_AWLEN[2] = hps2fpga_AWLEN_bus[2];
assign h2f_AWLEN[3] = hps2fpga_AWLEN_bus[3];

assign h2f_AWSIZE[0] = hps2fpga_AWSIZE_bus[0];
assign h2f_AWSIZE[1] = hps2fpga_AWSIZE_bus[1];
assign h2f_AWSIZE[2] = hps2fpga_AWSIZE_bus[2];

assign h2f_WDATA[0] = hps2fpga_WDATA_bus[0];
assign h2f_WDATA[1] = hps2fpga_WDATA_bus[1];
assign h2f_WDATA[2] = hps2fpga_WDATA_bus[2];
assign h2f_WDATA[3] = hps2fpga_WDATA_bus[3];
assign h2f_WDATA[4] = hps2fpga_WDATA_bus[4];
assign h2f_WDATA[5] = hps2fpga_WDATA_bus[5];
assign h2f_WDATA[6] = hps2fpga_WDATA_bus[6];
assign h2f_WDATA[7] = hps2fpga_WDATA_bus[7];
assign h2f_WDATA[8] = hps2fpga_WDATA_bus[8];
assign h2f_WDATA[9] = hps2fpga_WDATA_bus[9];
assign h2f_WDATA[10] = hps2fpga_WDATA_bus[10];
assign h2f_WDATA[11] = hps2fpga_WDATA_bus[11];
assign h2f_WDATA[12] = hps2fpga_WDATA_bus[12];
assign h2f_WDATA[13] = hps2fpga_WDATA_bus[13];
assign h2f_WDATA[14] = hps2fpga_WDATA_bus[14];
assign h2f_WDATA[15] = hps2fpga_WDATA_bus[15];
assign h2f_WDATA[16] = hps2fpga_WDATA_bus[16];
assign h2f_WDATA[17] = hps2fpga_WDATA_bus[17];
assign h2f_WDATA[18] = hps2fpga_WDATA_bus[18];
assign h2f_WDATA[19] = hps2fpga_WDATA_bus[19];
assign h2f_WDATA[20] = hps2fpga_WDATA_bus[20];
assign h2f_WDATA[21] = hps2fpga_WDATA_bus[21];
assign h2f_WDATA[22] = hps2fpga_WDATA_bus[22];
assign h2f_WDATA[23] = hps2fpga_WDATA_bus[23];
assign h2f_WDATA[24] = hps2fpga_WDATA_bus[24];
assign h2f_WDATA[25] = hps2fpga_WDATA_bus[25];
assign h2f_WDATA[26] = hps2fpga_WDATA_bus[26];
assign h2f_WDATA[27] = hps2fpga_WDATA_bus[27];
assign h2f_WDATA[28] = hps2fpga_WDATA_bus[28];
assign h2f_WDATA[29] = hps2fpga_WDATA_bus[29];
assign h2f_WDATA[30] = hps2fpga_WDATA_bus[30];
assign h2f_WDATA[31] = hps2fpga_WDATA_bus[31];
assign h2f_WDATA[32] = hps2fpga_WDATA_bus[32];
assign h2f_WDATA[33] = hps2fpga_WDATA_bus[33];
assign h2f_WDATA[34] = hps2fpga_WDATA_bus[34];
assign h2f_WDATA[35] = hps2fpga_WDATA_bus[35];
assign h2f_WDATA[36] = hps2fpga_WDATA_bus[36];
assign h2f_WDATA[37] = hps2fpga_WDATA_bus[37];
assign h2f_WDATA[38] = hps2fpga_WDATA_bus[38];
assign h2f_WDATA[39] = hps2fpga_WDATA_bus[39];
assign h2f_WDATA[40] = hps2fpga_WDATA_bus[40];
assign h2f_WDATA[41] = hps2fpga_WDATA_bus[41];
assign h2f_WDATA[42] = hps2fpga_WDATA_bus[42];
assign h2f_WDATA[43] = hps2fpga_WDATA_bus[43];
assign h2f_WDATA[44] = hps2fpga_WDATA_bus[44];
assign h2f_WDATA[45] = hps2fpga_WDATA_bus[45];
assign h2f_WDATA[46] = hps2fpga_WDATA_bus[46];
assign h2f_WDATA[47] = hps2fpga_WDATA_bus[47];
assign h2f_WDATA[48] = hps2fpga_WDATA_bus[48];
assign h2f_WDATA[49] = hps2fpga_WDATA_bus[49];
assign h2f_WDATA[50] = hps2fpga_WDATA_bus[50];
assign h2f_WDATA[51] = hps2fpga_WDATA_bus[51];
assign h2f_WDATA[52] = hps2fpga_WDATA_bus[52];
assign h2f_WDATA[53] = hps2fpga_WDATA_bus[53];
assign h2f_WDATA[54] = hps2fpga_WDATA_bus[54];
assign h2f_WDATA[55] = hps2fpga_WDATA_bus[55];
assign h2f_WDATA[56] = hps2fpga_WDATA_bus[56];
assign h2f_WDATA[57] = hps2fpga_WDATA_bus[57];
assign h2f_WDATA[58] = hps2fpga_WDATA_bus[58];
assign h2f_WDATA[59] = hps2fpga_WDATA_bus[59];
assign h2f_WDATA[60] = hps2fpga_WDATA_bus[60];
assign h2f_WDATA[61] = hps2fpga_WDATA_bus[61];
assign h2f_WDATA[62] = hps2fpga_WDATA_bus[62];
assign h2f_WDATA[63] = hps2fpga_WDATA_bus[63];
assign h2f_WDATA[64] = hps2fpga_WDATA_bus[64];
assign h2f_WDATA[65] = hps2fpga_WDATA_bus[65];
assign h2f_WDATA[66] = hps2fpga_WDATA_bus[66];
assign h2f_WDATA[67] = hps2fpga_WDATA_bus[67];
assign h2f_WDATA[68] = hps2fpga_WDATA_bus[68];
assign h2f_WDATA[69] = hps2fpga_WDATA_bus[69];
assign h2f_WDATA[70] = hps2fpga_WDATA_bus[70];
assign h2f_WDATA[71] = hps2fpga_WDATA_bus[71];
assign h2f_WDATA[72] = hps2fpga_WDATA_bus[72];
assign h2f_WDATA[73] = hps2fpga_WDATA_bus[73];
assign h2f_WDATA[74] = hps2fpga_WDATA_bus[74];
assign h2f_WDATA[75] = hps2fpga_WDATA_bus[75];
assign h2f_WDATA[76] = hps2fpga_WDATA_bus[76];
assign h2f_WDATA[77] = hps2fpga_WDATA_bus[77];
assign h2f_WDATA[78] = hps2fpga_WDATA_bus[78];
assign h2f_WDATA[79] = hps2fpga_WDATA_bus[79];
assign h2f_WDATA[80] = hps2fpga_WDATA_bus[80];
assign h2f_WDATA[81] = hps2fpga_WDATA_bus[81];
assign h2f_WDATA[82] = hps2fpga_WDATA_bus[82];
assign h2f_WDATA[83] = hps2fpga_WDATA_bus[83];
assign h2f_WDATA[84] = hps2fpga_WDATA_bus[84];
assign h2f_WDATA[85] = hps2fpga_WDATA_bus[85];
assign h2f_WDATA[86] = hps2fpga_WDATA_bus[86];
assign h2f_WDATA[87] = hps2fpga_WDATA_bus[87];
assign h2f_WDATA[88] = hps2fpga_WDATA_bus[88];
assign h2f_WDATA[89] = hps2fpga_WDATA_bus[89];
assign h2f_WDATA[90] = hps2fpga_WDATA_bus[90];
assign h2f_WDATA[91] = hps2fpga_WDATA_bus[91];
assign h2f_WDATA[92] = hps2fpga_WDATA_bus[92];
assign h2f_WDATA[93] = hps2fpga_WDATA_bus[93];
assign h2f_WDATA[94] = hps2fpga_WDATA_bus[94];
assign h2f_WDATA[95] = hps2fpga_WDATA_bus[95];
assign h2f_WDATA[96] = hps2fpga_WDATA_bus[96];
assign h2f_WDATA[97] = hps2fpga_WDATA_bus[97];
assign h2f_WDATA[98] = hps2fpga_WDATA_bus[98];
assign h2f_WDATA[99] = hps2fpga_WDATA_bus[99];
assign h2f_WDATA[100] = hps2fpga_WDATA_bus[100];
assign h2f_WDATA[101] = hps2fpga_WDATA_bus[101];
assign h2f_WDATA[102] = hps2fpga_WDATA_bus[102];
assign h2f_WDATA[103] = hps2fpga_WDATA_bus[103];
assign h2f_WDATA[104] = hps2fpga_WDATA_bus[104];
assign h2f_WDATA[105] = hps2fpga_WDATA_bus[105];
assign h2f_WDATA[106] = hps2fpga_WDATA_bus[106];
assign h2f_WDATA[107] = hps2fpga_WDATA_bus[107];
assign h2f_WDATA[108] = hps2fpga_WDATA_bus[108];
assign h2f_WDATA[109] = hps2fpga_WDATA_bus[109];
assign h2f_WDATA[110] = hps2fpga_WDATA_bus[110];
assign h2f_WDATA[111] = hps2fpga_WDATA_bus[111];
assign h2f_WDATA[112] = hps2fpga_WDATA_bus[112];
assign h2f_WDATA[113] = hps2fpga_WDATA_bus[113];
assign h2f_WDATA[114] = hps2fpga_WDATA_bus[114];
assign h2f_WDATA[115] = hps2fpga_WDATA_bus[115];
assign h2f_WDATA[116] = hps2fpga_WDATA_bus[116];
assign h2f_WDATA[117] = hps2fpga_WDATA_bus[117];
assign h2f_WDATA[118] = hps2fpga_WDATA_bus[118];
assign h2f_WDATA[119] = hps2fpga_WDATA_bus[119];
assign h2f_WDATA[120] = hps2fpga_WDATA_bus[120];
assign h2f_WDATA[121] = hps2fpga_WDATA_bus[121];
assign h2f_WDATA[122] = hps2fpga_WDATA_bus[122];
assign h2f_WDATA[123] = hps2fpga_WDATA_bus[123];
assign h2f_WDATA[124] = hps2fpga_WDATA_bus[124];
assign h2f_WDATA[125] = hps2fpga_WDATA_bus[125];
assign h2f_WDATA[126] = hps2fpga_WDATA_bus[126];
assign h2f_WDATA[127] = hps2fpga_WDATA_bus[127];

assign h2f_WSTRB[0] = hps2fpga_WSTRB_bus[0];
assign h2f_WSTRB[1] = hps2fpga_WSTRB_bus[1];
assign h2f_WSTRB[2] = hps2fpga_WSTRB_bus[2];
assign h2f_WSTRB[3] = hps2fpga_WSTRB_bus[3];
assign h2f_WSTRB[4] = hps2fpga_WSTRB_bus[4];
assign h2f_WSTRB[5] = hps2fpga_WSTRB_bus[5];
assign h2f_WSTRB[6] = hps2fpga_WSTRB_bus[6];
assign h2f_WSTRB[7] = hps2fpga_WSTRB_bus[7];
assign h2f_WSTRB[8] = hps2fpga_WSTRB_bus[8];
assign h2f_WSTRB[9] = hps2fpga_WSTRB_bus[9];
assign h2f_WSTRB[10] = hps2fpga_WSTRB_bus[10];
assign h2f_WSTRB[11] = hps2fpga_WSTRB_bus[11];
assign h2f_WSTRB[12] = hps2fpga_WSTRB_bus[12];
assign h2f_WSTRB[13] = hps2fpga_WSTRB_bus[13];
assign h2f_WSTRB[14] = hps2fpga_WSTRB_bus[14];
assign h2f_WSTRB[15] = hps2fpga_WSTRB_bus[15];

cyclonev_hps_interface_clocks_resets clocks_resets(
	.f2h_cold_rst_req_n(vcc),
	.f2h_dbg_rst_req_n(vcc),
	.f2h_pending_rst_ack(vcc),
	.f2h_periph_ref_clk(gnd),
	.f2h_sdram_ref_clk(gnd),
	.f2h_warm_rst_req_n(vcc),
	.ptp_ref_clk(gnd),
	.h2f_cold_rst_n(\clocks_resets~h2f_cold_rst_n ),
	.h2f_pending_rst_req_n(),
	.h2f_rst_n(h2f_rst_n[0]),
	.h2f_user0_clk(),
	.h2f_user1_clk(),
	.h2f_user2_clk());
defparam clocks_resets.h2f_user0_clk_freq = 100;
defparam clocks_resets.h2f_user1_clk_freq = 100;
defparam clocks_resets.h2f_user2_clk_freq = 100;

cyclonev_hps_interface_hps2fpga_light_weight hps2fpga_light_weight(
	.arready(h2f_lw_ARREADY[0]),
	.awready(h2f_lw_AWREADY[0]),
	.bvalid(h2f_lw_BVALID[0]),
	.clk(h2f_lw_axi_clk[0]),
	.rlast(h2f_lw_RLAST[0]),
	.rvalid(h2f_lw_RVALID[0]),
	.wready(h2f_lw_WREADY[0]),
	.bid({h2f_lw_BID[11],h2f_lw_BID[10],h2f_lw_BID[9],h2f_lw_BID[8],h2f_lw_BID[7],h2f_lw_BID[6],h2f_lw_BID[5],h2f_lw_BID[4],h2f_lw_BID[3],h2f_lw_BID[2],h2f_lw_BID[1],h2f_lw_BID[0]}),
	.bresp({gnd,gnd}),
	.rdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,h2f_lw_RDATA[7],h2f_lw_RDATA[6],h2f_lw_RDATA[5],h2f_lw_RDATA[4],h2f_lw_RDATA[3],h2f_lw_RDATA[2],h2f_lw_RDATA[1],h2f_lw_RDATA[0]}),
	.rid({h2f_lw_BID[11],h2f_lw_BID[10],h2f_lw_BID[9],h2f_lw_BID[8],h2f_lw_BID[7],h2f_lw_BID[6],h2f_lw_BID[5],h2f_lw_BID[4],h2f_lw_BID[3],h2f_lw_BID[2],h2f_lw_BID[1],h2f_lw_BID[0]}),
	.rresp({gnd,gnd}),
	.arvalid(h2f_lw_ARVALID[0]),
	.awvalid(h2f_lw_AWVALID[0]),
	.bready(h2f_lw_BREADY[0]),
	.rready(h2f_lw_RREADY[0]),
	.wlast(h2f_lw_WLAST[0]),
	.wvalid(h2f_lw_WVALID[0]),
	.araddr(hps2fpga_light_weight_ARADDR_bus),
	.arburst(hps2fpga_light_weight_ARBURST_bus),
	.arcache(),
	.arid(hps2fpga_light_weight_ARID_bus),
	.arlen(hps2fpga_light_weight_ARLEN_bus),
	.arlock(),
	.arprot(),
	.arsize(hps2fpga_light_weight_ARSIZE_bus),
	.awaddr(hps2fpga_light_weight_AWADDR_bus),
	.awburst(hps2fpga_light_weight_AWBURST_bus),
	.awcache(),
	.awid(hps2fpga_light_weight_AWID_bus),
	.awlen(hps2fpga_light_weight_AWLEN_bus),
	.awlock(),
	.awprot(),
	.awsize(hps2fpga_light_weight_AWSIZE_bus),
	.wdata(hps2fpga_light_weight_WDATA_bus),
	.wid(),
	.wstrb(hps2fpga_light_weight_WSTRB_bus));

cyclonev_hps_interface_hps2fpga hps2fpga(
	.arready(h2f_ARREADY[0]),
	.awready(h2f_AWREADY[0]),
	.bvalid(h2f_BVALID[0]),
	.clk(h2f_lw_axi_clk[0]),
	.rlast(h2f_RLAST[0]),
	.rvalid(h2f_RVALID[0]),
	.wready(h2f_WREADY[0]),
	.bid({h2f_BID[11],h2f_BID[10],h2f_BID[9],h2f_BID[8],h2f_BID[7],h2f_BID[6],h2f_BID[5],h2f_BID[4],h2f_BID[3],h2f_BID[2],h2f_BID[1],h2f_BID[0]}),
	.bresp({gnd,gnd}),
	.port_size_config({vcc,gnd}),
	.rdata({h2f_RDATA[127],h2f_RDATA[126],h2f_RDATA[125],h2f_RDATA[124],h2f_RDATA[123],h2f_RDATA[122],h2f_RDATA[121],h2f_RDATA[120],h2f_RDATA[119],h2f_RDATA[118],h2f_RDATA[117],h2f_RDATA[116],h2f_RDATA[115],h2f_RDATA[114],h2f_RDATA[113],h2f_RDATA[112],h2f_RDATA[111],h2f_RDATA[110],h2f_RDATA[109],h2f_RDATA[108],h2f_RDATA[107],h2f_RDATA[106],h2f_RDATA[105],h2f_RDATA[104],h2f_RDATA[103],h2f_RDATA[102],h2f_RDATA[101],h2f_RDATA[100],
h2f_RDATA[99],h2f_RDATA[98],h2f_RDATA[97],h2f_RDATA[96],h2f_RDATA[95],h2f_RDATA[94],h2f_RDATA[93],h2f_RDATA[92],h2f_RDATA[91],h2f_RDATA[90],h2f_RDATA[89],h2f_RDATA[88],h2f_RDATA[87],h2f_RDATA[86],h2f_RDATA[85],h2f_RDATA[84],h2f_RDATA[83],h2f_RDATA[82],h2f_RDATA[81],h2f_RDATA[80],h2f_RDATA[79],h2f_RDATA[78],h2f_RDATA[77],h2f_RDATA[76],h2f_RDATA[75],h2f_RDATA[74],h2f_RDATA[73],h2f_RDATA[72],
h2f_RDATA[71],h2f_RDATA[70],h2f_RDATA[69],h2f_RDATA[68],h2f_RDATA[67],h2f_RDATA[66],h2f_RDATA[65],h2f_RDATA[64],h2f_RDATA[63],h2f_RDATA[62],h2f_RDATA[61],h2f_RDATA[60],h2f_RDATA[59],h2f_RDATA[58],h2f_RDATA[57],h2f_RDATA[56],h2f_RDATA[55],h2f_RDATA[54],h2f_RDATA[53],h2f_RDATA[52],h2f_RDATA[51],h2f_RDATA[50],h2f_RDATA[49],h2f_RDATA[48],h2f_RDATA[47],h2f_RDATA[46],h2f_RDATA[45],h2f_RDATA[44],
h2f_RDATA[43],h2f_RDATA[42],h2f_RDATA[41],h2f_RDATA[40],h2f_RDATA[39],h2f_RDATA[38],h2f_RDATA[37],h2f_RDATA[36],h2f_RDATA[35],h2f_RDATA[34],h2f_RDATA[33],h2f_RDATA[32],h2f_RDATA[31],h2f_RDATA[30],h2f_RDATA[29],h2f_RDATA[28],h2f_RDATA[27],h2f_RDATA[26],h2f_RDATA[25],h2f_RDATA[24],h2f_RDATA[23],h2f_RDATA[22],h2f_RDATA[21],h2f_RDATA[20],h2f_RDATA[19],h2f_RDATA[18],h2f_RDATA[17],h2f_RDATA[16],
h2f_RDATA[15],h2f_RDATA[14],h2f_RDATA[13],h2f_RDATA[12],h2f_RDATA[11],h2f_RDATA[10],h2f_RDATA[9],h2f_RDATA[8],h2f_RDATA[7],h2f_RDATA[6],h2f_RDATA[5],h2f_RDATA[4],h2f_RDATA[3],h2f_RDATA[2],h2f_RDATA[1],h2f_RDATA[0]}),
	.rid({h2f_RID[11],h2f_RID[10],h2f_RID[9],h2f_RID[8],h2f_RID[7],h2f_RID[6],h2f_RID[5],h2f_RID[4],h2f_RID[3],h2f_RID[2],h2f_RID[1],h2f_RID[0]}),
	.rresp({gnd,gnd}),
	.arvalid(h2f_ARVALID[0]),
	.awvalid(h2f_AWVALID[0]),
	.bready(h2f_BREADY[0]),
	.rready(h2f_RREADY[0]),
	.wlast(h2f_WLAST[0]),
	.wvalid(h2f_WVALID[0]),
	.araddr(hps2fpga_ARADDR_bus),
	.arburst(hps2fpga_ARBURST_bus),
	.arcache(),
	.arid(hps2fpga_ARID_bus),
	.arlen(hps2fpga_ARLEN_bus),
	.arlock(),
	.arprot(),
	.arsize(hps2fpga_ARSIZE_bus),
	.awaddr(hps2fpga_AWADDR_bus),
	.awburst(hps2fpga_AWBURST_bus),
	.awcache(),
	.awid(hps2fpga_AWID_bus),
	.awlen(hps2fpga_AWLEN_bus),
	.awlock(),
	.awprot(),
	.awsize(hps2fpga_AWSIZE_bus),
	.wdata(hps2fpga_WDATA_bus),
	.wid(),
	.wstrb(hps2fpga_WSTRB_bus));
defparam hps2fpga.data_width = 32;

cyclonev_hps_interface_dbg_apb debug_apb(
	.p_slv_err(gnd),
	.p_ready(gnd),
	.p_clk(gnd),
	.p_clk_en(gnd),
	.dbg_apb_disable(gnd),
	.p_rdata(32'b00000000000000000000000000000000),
	.p_addr_31(\debug_apb~O_P_ADDR_31 ),
	.p_write(),
	.p_sel(),
	.p_enable(),
	.p_reset_n(),
	.p_addr(),
	.p_wdata());
defparam debug_apb.dummy_param = 256;

cyclonev_hps_interface_tpiu_trace tpiu(
	.traceclk_ctl(vcc),
	.traceclkin(gnd),
	.traceclk(),
	.trace_data(tpiu_TRACE_DATA_bus));

cyclonev_hps_interface_boot_from_fpga boot_from_fpga(
	.boot_from_fpga_on_failure(gnd),
	.boot_from_fpga_ready(gnd),
	.bsel_en(gnd),
	.csel_en(gnd),
	.bsel({gnd,gnd,vcc}),
	.csel({gnd,vcc}),
	.fake_dout(\boot_from_fpga~fake_dout ));

cyclonev_hps_interface_fpga2hps fpga2hps(
	.arvalid(gnd),
	.awvalid(gnd),
	.bready(gnd),
	.clk(h2f_lw_axi_clk[0]),
	.rready(gnd),
	.wlast(gnd),
	.wvalid(gnd),
	.araddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.arburst({gnd,gnd}),
	.arcache({gnd,gnd,gnd,gnd}),
	.arid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.arlen({gnd,gnd,gnd,gnd}),
	.arlock({gnd,gnd}),
	.arprot({gnd,gnd,gnd}),
	.arsize({gnd,gnd,gnd}),
	.aruser({gnd,gnd,gnd,gnd,gnd}),
	.awaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.awburst({gnd,gnd}),
	.awcache({gnd,gnd,gnd,gnd}),
	.awid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.awlen({gnd,gnd,gnd,gnd}),
	.awlock({gnd,gnd}),
	.awprot({gnd,gnd,gnd}),
	.awsize({gnd,gnd,gnd}),
	.awuser({gnd,gnd,gnd,gnd,gnd}),
	.port_size_config({gnd,vcc}),
	.wdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.wid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.wstrb({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.arready(\f2h_ARREADY[0] ),
	.awready(),
	.bvalid(),
	.rlast(),
	.rvalid(),
	.wready(),
	.bid(),
	.bresp(),
	.rdata(),
	.rid(),
	.rresp());
defparam fpga2hps.data_width = 32;

cyclonev_hps_interface_fpga2sdram f2sdram(
	.cmd_port_clk_0(gnd),
	.cmd_port_clk_1(gnd),
	.cmd_port_clk_2(gnd),
	.cmd_port_clk_3(gnd),
	.cmd_port_clk_4(gnd),
	.cmd_port_clk_5(gnd),
	.cmd_valid_0(gnd),
	.cmd_valid_1(gnd),
	.cmd_valid_2(gnd),
	.cmd_valid_3(gnd),
	.cmd_valid_4(gnd),
	.cmd_valid_5(gnd),
	.rd_clk_0(gnd),
	.rd_clk_1(gnd),
	.rd_clk_2(gnd),
	.rd_clk_3(gnd),
	.rd_ready_0(gnd),
	.rd_ready_1(gnd),
	.rd_ready_2(gnd),
	.rd_ready_3(gnd),
	.wr_clk_0(gnd),
	.wr_clk_1(gnd),
	.wr_clk_2(gnd),
	.wr_clk_3(gnd),
	.wr_valid_0(gnd),
	.wr_valid_1(gnd),
	.wr_valid_2(gnd),
	.wr_valid_3(gnd),
	.wrack_ready_0(gnd),
	.wrack_ready_1(gnd),
	.wrack_ready_2(gnd),
	.wrack_ready_3(gnd),
	.wrack_ready_4(gnd),
	.wrack_ready_5(gnd),
	.cfg_axi_mm_select({gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_rfifo_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_type({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_wfifo_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_port_width({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_rfifo_cport_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_wfifo_cport_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cmd_data_0(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_1(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_2(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_3(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_4(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_5(60'b000000000000000000000000000000000000000000000000000000000000),
	.wr_data_0(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_1(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_2(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.wr_data_3(90'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
	.cmd_ready_0(),
	.cmd_ready_1(),
	.cmd_ready_2(),
	.cmd_ready_3(),
	.cmd_ready_4(),
	.cmd_ready_5(),
	.rd_valid_0(),
	.rd_valid_1(),
	.rd_valid_2(),
	.rd_valid_3(),
	.wr_ready_0(),
	.wr_ready_1(),
	.wr_ready_2(),
	.wr_ready_3(),
	.wrack_valid_0(),
	.wrack_valid_1(),
	.wrack_valid_2(),
	.wrack_valid_3(),
	.wrack_valid_4(),
	.wrack_valid_5(),
	.bonding_out_1(f2sdram_BONDING_OUT_1_bus),
	.bonding_out_2(),
	.rd_data_0(),
	.rd_data_1(),
	.rd_data_2(),
	.rd_data_3(),
	.wrack_data_0(),
	.wrack_data_1(),
	.wrack_data_2(),
	.wrack_data_3(),
	.wrack_data_4(),
	.wrack_data_5());

cyclonev_hps_interface_interrupts interrupts(
	.irq({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.fake_dout(\interrupts~fake_dout ),
	.h2f_can0_irq(),
	.h2f_can1_irq(),
	.h2f_clkmgr_irq(),
	.h2f_cti_irq0_n(),
	.h2f_cti_irq1_n(),
	.h2f_dma_abort_irq(),
	.h2f_dma_irq0(),
	.h2f_dma_irq1(),
	.h2f_dma_irq2(),
	.h2f_dma_irq3(),
	.h2f_dma_irq4(),
	.h2f_dma_irq5(),
	.h2f_dma_irq6(),
	.h2f_dma_irq7(),
	.h2f_emac0_irq(),
	.h2f_emac1_irq(),
	.h2f_fpga_man_irq(),
	.h2f_gpio0_irq(),
	.h2f_gpio1_irq(),
	.h2f_gpio2_irq(),
	.h2f_i2c0_irq(),
	.h2f_i2c1_irq(),
	.h2f_i2c_emac0_irq(),
	.h2f_i2c_emac1_irq(),
	.h2f_l4sp0_irq(),
	.h2f_l4sp1_irq(),
	.h2f_mpuwakeup_irq(),
	.h2f_nand_irq(),
	.h2f_osc0_irq(),
	.h2f_osc1_irq(),
	.h2f_qspi_irq(),
	.h2f_sdmmc_irq(),
	.h2f_spi0_irq(),
	.h2f_spi1_irq(),
	.h2f_spi2_irq(),
	.h2f_spi3_irq(),
	.h2f_uart0_irq(),
	.h2f_uart1_irq(),
	.h2f_usb0_irq(),
	.h2f_usb1_irq(),
	.h2f_wdog0_irq(),
	.h2f_wdog1_irq());

endmodule

module Computer_System_Computer_System_ARM_A9_HPS_hps_io (
	emac1_inst,
	emac1_inst1,
	intermediate_0,
	intermediate_1,
	emac1_inst2,
	emac1_inst3,
	emac1_inst4,
	emac1_inst5,
	emac1_inst6,
	qspi_inst,
	intermediate_2,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_3,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	qspi_inst1,
	sdio_inst,
	intermediate_10,
	intermediate_11,
	intermediate_12,
	intermediate_14,
	intermediate_16,
	intermediate_18,
	intermediate_13,
	intermediate_15,
	intermediate_17,
	intermediate_19,
	usb1_inst,
	intermediate_20,
	intermediate_22,
	intermediate_24,
	intermediate_26,
	intermediate_28,
	intermediate_30,
	intermediate_32,
	intermediate_34,
	intermediate_21,
	intermediate_23,
	intermediate_25,
	intermediate_27,
	intermediate_29,
	intermediate_31,
	intermediate_33,
	intermediate_35,
	spim1_inst,
	spim1_inst1,
	intermediate_36,
	intermediate_37,
	uart0_inst,
	intermediate_39,
	intermediate_38,
	intermediate_41,
	intermediate_40,
	intermediate_42,
	intermediate_43,
	intermediate_44,
	intermediate_46,
	intermediate_48,
	intermediate_50,
	intermediate_52,
	intermediate_54,
	intermediate_45,
	intermediate_47,
	intermediate_49,
	intermediate_51,
	intermediate_53,
	intermediate_55,
	intermediate_56,
	intermediate_57,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_qspi_inst_IO0_0,
	hps_io_qspi_inst_IO1_0,
	hps_io_qspi_inst_IO2_0,
	hps_io_qspi_inst_IO3_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_io_usb1_inst_D0_0,
	hps_io_usb1_inst_D1_0,
	hps_io_usb1_inst_D2_0,
	hps_io_usb1_inst_D3_0,
	hps_io_usb1_inst_D4_0,
	hps_io_usb1_inst_D5_0,
	hps_io_usb1_inst_D6_0,
	hps_io_usb1_inst_D7_0,
	hps_io_i2c0_inst_SDA_0,
	hps_io_i2c0_inst_SCL_0,
	hps_io_i2c1_inst_SDA_0,
	hps_io_i2c1_inst_SCL_0,
	hps_io_gpio_inst_GPIO09_0,
	hps_io_gpio_inst_GPIO35_0,
	hps_io_gpio_inst_GPIO40_0,
	hps_io_gpio_inst_GPIO41_0,
	hps_io_gpio_inst_GPIO48_0,
	hps_io_gpio_inst_GPIO53_0,
	hps_io_gpio_inst_GPIO54_0,
	hps_io_gpio_inst_GPIO61_0,
	hps_io_hps_io_emac1_inst_RXD0,
	hps_io_hps_io_emac1_inst_RXD1,
	hps_io_hps_io_emac1_inst_RXD2,
	hps_io_hps_io_emac1_inst_RXD3,
	hps_io_hps_io_emac1_inst_RX_CLK,
	hps_io_hps_io_emac1_inst_RX_CTL,
	hps_io_hps_io_spim1_inst_MISO,
	hps_io_hps_io_uart0_inst_RX,
	hps_io_hps_io_usb1_inst_CLK,
	hps_io_hps_io_usb1_inst_DIR,
	hps_io_hps_io_usb1_inst_NXT,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	emac1_inst;
output 	emac1_inst1;
output 	intermediate_0;
output 	intermediate_1;
output 	emac1_inst2;
output 	emac1_inst3;
output 	emac1_inst4;
output 	emac1_inst5;
output 	emac1_inst6;
output 	qspi_inst;
output 	intermediate_2;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_3;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	qspi_inst1;
output 	sdio_inst;
output 	intermediate_10;
output 	intermediate_11;
output 	intermediate_12;
output 	intermediate_14;
output 	intermediate_16;
output 	intermediate_18;
output 	intermediate_13;
output 	intermediate_15;
output 	intermediate_17;
output 	intermediate_19;
output 	usb1_inst;
output 	intermediate_20;
output 	intermediate_22;
output 	intermediate_24;
output 	intermediate_26;
output 	intermediate_28;
output 	intermediate_30;
output 	intermediate_32;
output 	intermediate_34;
output 	intermediate_21;
output 	intermediate_23;
output 	intermediate_25;
output 	intermediate_27;
output 	intermediate_29;
output 	intermediate_31;
output 	intermediate_33;
output 	intermediate_35;
output 	spim1_inst;
output 	spim1_inst1;
output 	intermediate_36;
output 	intermediate_37;
output 	uart0_inst;
output 	intermediate_39;
output 	intermediate_38;
output 	intermediate_41;
output 	intermediate_40;
output 	intermediate_42;
output 	intermediate_43;
output 	intermediate_44;
output 	intermediate_46;
output 	intermediate_48;
output 	intermediate_50;
output 	intermediate_52;
output 	intermediate_54;
output 	intermediate_45;
output 	intermediate_47;
output 	intermediate_49;
output 	intermediate_51;
output 	intermediate_53;
output 	intermediate_55;
output 	intermediate_56;
output 	intermediate_57;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_qspi_inst_IO0_0;
input 	hps_io_qspi_inst_IO1_0;
input 	hps_io_qspi_inst_IO2_0;
input 	hps_io_qspi_inst_IO3_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_io_usb1_inst_D0_0;
input 	hps_io_usb1_inst_D1_0;
input 	hps_io_usb1_inst_D2_0;
input 	hps_io_usb1_inst_D3_0;
input 	hps_io_usb1_inst_D4_0;
input 	hps_io_usb1_inst_D5_0;
input 	hps_io_usb1_inst_D6_0;
input 	hps_io_usb1_inst_D7_0;
input 	hps_io_i2c0_inst_SDA_0;
input 	hps_io_i2c0_inst_SCL_0;
input 	hps_io_i2c1_inst_SDA_0;
input 	hps_io_i2c1_inst_SCL_0;
input 	hps_io_gpio_inst_GPIO09_0;
input 	hps_io_gpio_inst_GPIO35_0;
input 	hps_io_gpio_inst_GPIO40_0;
input 	hps_io_gpio_inst_GPIO41_0;
input 	hps_io_gpio_inst_GPIO48_0;
input 	hps_io_gpio_inst_GPIO53_0;
input 	hps_io_gpio_inst_GPIO54_0;
input 	hps_io_gpio_inst_GPIO61_0;
input 	hps_io_hps_io_emac1_inst_RXD0;
input 	hps_io_hps_io_emac1_inst_RXD1;
input 	hps_io_hps_io_emac1_inst_RXD2;
input 	hps_io_hps_io_emac1_inst_RXD3;
input 	hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_io_hps_io_emac1_inst_RX_CTL;
input 	hps_io_hps_io_spim1_inst_MISO;
input 	hps_io_hps_io_uart0_inst_RX;
input 	hps_io_hps_io_usb1_inst_CLK;
input 	hps_io_hps_io_usb1_inst_DIR;
input 	hps_io_hps_io_usb1_inst_NXT;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_Computer_System_ARM_A9_HPS_hps_io_border border(
	.hps_io_emac1_inst_TX_CLK({emac1_inst}),
	.hps_io_emac1_inst_TX_CTL({emac1_inst1}),
	.intermediate_0(intermediate_0),
	.intermediate_1(intermediate_1),
	.hps_io_emac1_inst_MDC({emac1_inst2}),
	.hps_io_emac1_inst_TXD0({emac1_inst3}),
	.hps_io_emac1_inst_TXD1({emac1_inst4}),
	.hps_io_emac1_inst_TXD2({emac1_inst5}),
	.hps_io_emac1_inst_TXD3({emac1_inst6}),
	.hps_io_qspi_inst_CLK({qspi_inst}),
	.intermediate_2(intermediate_2),
	.intermediate_4(intermediate_4),
	.intermediate_6(intermediate_6),
	.intermediate_8(intermediate_8),
	.intermediate_3(intermediate_3),
	.intermediate_5(intermediate_5),
	.intermediate_7(intermediate_7),
	.intermediate_9(intermediate_9),
	.hps_io_qspi_inst_SS0({qspi_inst1}),
	.hps_io_sdio_inst_CLK({sdio_inst}),
	.intermediate_10(intermediate_10),
	.intermediate_11(intermediate_11),
	.intermediate_12(intermediate_12),
	.intermediate_14(intermediate_14),
	.intermediate_16(intermediate_16),
	.intermediate_18(intermediate_18),
	.intermediate_13(intermediate_13),
	.intermediate_15(intermediate_15),
	.intermediate_17(intermediate_17),
	.intermediate_19(intermediate_19),
	.hps_io_usb1_inst_STP({usb1_inst}),
	.intermediate_20(intermediate_20),
	.intermediate_22(intermediate_22),
	.intermediate_24(intermediate_24),
	.intermediate_26(intermediate_26),
	.intermediate_28(intermediate_28),
	.intermediate_30(intermediate_30),
	.intermediate_32(intermediate_32),
	.intermediate_34(intermediate_34),
	.intermediate_21(intermediate_21),
	.intermediate_23(intermediate_23),
	.intermediate_25(intermediate_25),
	.intermediate_27(intermediate_27),
	.intermediate_29(intermediate_29),
	.intermediate_31(intermediate_31),
	.intermediate_33(intermediate_33),
	.intermediate_35(intermediate_35),
	.hps_io_spim1_inst_CLK({spim1_inst}),
	.hps_io_spim1_inst_SS0({spim1_inst1}),
	.intermediate_36(intermediate_36),
	.intermediate_37(intermediate_37),
	.hps_io_uart0_inst_TX({uart0_inst}),
	.intermediate_39(intermediate_39),
	.intermediate_38(intermediate_38),
	.intermediate_41(intermediate_41),
	.intermediate_40(intermediate_40),
	.intermediate_42(intermediate_42),
	.intermediate_43(intermediate_43),
	.intermediate_44(intermediate_44),
	.intermediate_46(intermediate_46),
	.intermediate_48(intermediate_48),
	.intermediate_50(intermediate_50),
	.intermediate_52(intermediate_52),
	.intermediate_54(intermediate_54),
	.intermediate_45(intermediate_45),
	.intermediate_47(intermediate_47),
	.intermediate_49(intermediate_49),
	.intermediate_51(intermediate_51),
	.intermediate_53(intermediate_53),
	.intermediate_55(intermediate_55),
	.intermediate_56(intermediate_56),
	.intermediate_57(intermediate_57),
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.hps_io_emac1_inst_MDIO_0(hps_io_emac1_inst_MDIO_0),
	.hps_io_qspi_inst_IO0_0(hps_io_qspi_inst_IO0_0),
	.hps_io_qspi_inst_IO1_0(hps_io_qspi_inst_IO1_0),
	.hps_io_qspi_inst_IO2_0(hps_io_qspi_inst_IO2_0),
	.hps_io_qspi_inst_IO3_0(hps_io_qspi_inst_IO3_0),
	.hps_io_sdio_inst_CMD_0(hps_io_sdio_inst_CMD_0),
	.hps_io_sdio_inst_D0_0(hps_io_sdio_inst_D0_0),
	.hps_io_sdio_inst_D1_0(hps_io_sdio_inst_D1_0),
	.hps_io_sdio_inst_D2_0(hps_io_sdio_inst_D2_0),
	.hps_io_sdio_inst_D3_0(hps_io_sdio_inst_D3_0),
	.hps_io_usb1_inst_D0_0(hps_io_usb1_inst_D0_0),
	.hps_io_usb1_inst_D1_0(hps_io_usb1_inst_D1_0),
	.hps_io_usb1_inst_D2_0(hps_io_usb1_inst_D2_0),
	.hps_io_usb1_inst_D3_0(hps_io_usb1_inst_D3_0),
	.hps_io_usb1_inst_D4_0(hps_io_usb1_inst_D4_0),
	.hps_io_usb1_inst_D5_0(hps_io_usb1_inst_D5_0),
	.hps_io_usb1_inst_D6_0(hps_io_usb1_inst_D6_0),
	.hps_io_usb1_inst_D7_0(hps_io_usb1_inst_D7_0),
	.hps_io_i2c0_inst_SDA_0(hps_io_i2c0_inst_SDA_0),
	.hps_io_i2c0_inst_SCL_0(hps_io_i2c0_inst_SCL_0),
	.hps_io_i2c1_inst_SDA_0(hps_io_i2c1_inst_SDA_0),
	.hps_io_i2c1_inst_SCL_0(hps_io_i2c1_inst_SCL_0),
	.hps_io_gpio_inst_GPIO09_0(hps_io_gpio_inst_GPIO09_0),
	.hps_io_gpio_inst_GPIO35_0(hps_io_gpio_inst_GPIO35_0),
	.hps_io_gpio_inst_GPIO40_0(hps_io_gpio_inst_GPIO40_0),
	.hps_io_gpio_inst_GPIO41_0(hps_io_gpio_inst_GPIO41_0),
	.hps_io_gpio_inst_GPIO48_0(hps_io_gpio_inst_GPIO48_0),
	.hps_io_gpio_inst_GPIO53_0(hps_io_gpio_inst_GPIO53_0),
	.hps_io_gpio_inst_GPIO54_0(hps_io_gpio_inst_GPIO54_0),
	.hps_io_gpio_inst_GPIO61_0(hps_io_gpio_inst_GPIO61_0),
	.hps_io_emac1_inst_RXD0({hps_io_hps_io_emac1_inst_RXD0}),
	.hps_io_emac1_inst_RXD1({hps_io_hps_io_emac1_inst_RXD1}),
	.hps_io_emac1_inst_RXD2({hps_io_hps_io_emac1_inst_RXD2}),
	.hps_io_emac1_inst_RXD3({hps_io_hps_io_emac1_inst_RXD3}),
	.hps_io_emac1_inst_RX_CLK({hps_io_hps_io_emac1_inst_RX_CLK}),
	.hps_io_emac1_inst_RX_CTL({hps_io_hps_io_emac1_inst_RX_CTL}),
	.hps_io_spim1_inst_MISO({hps_io_hps_io_spim1_inst_MISO}),
	.hps_io_uart0_inst_RX({hps_io_hps_io_uart0_inst_RX}),
	.hps_io_usb1_inst_CLK({hps_io_hps_io_usb1_inst_CLK}),
	.hps_io_usb1_inst_DIR({hps_io_hps_io_usb1_inst_DIR}),
	.hps_io_usb1_inst_NXT({hps_io_hps_io_usb1_inst_NXT}),
	.memory_oct_rzqin(memory_oct_rzqin));

endmodule

module Computer_System_Computer_System_ARM_A9_HPS_hps_io_border (
	hps_io_emac1_inst_TX_CLK,
	hps_io_emac1_inst_TX_CTL,
	intermediate_0,
	intermediate_1,
	hps_io_emac1_inst_MDC,
	hps_io_emac1_inst_TXD0,
	hps_io_emac1_inst_TXD1,
	hps_io_emac1_inst_TXD2,
	hps_io_emac1_inst_TXD3,
	hps_io_qspi_inst_CLK,
	intermediate_2,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_3,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	hps_io_qspi_inst_SS0,
	hps_io_sdio_inst_CLK,
	intermediate_10,
	intermediate_11,
	intermediate_12,
	intermediate_14,
	intermediate_16,
	intermediate_18,
	intermediate_13,
	intermediate_15,
	intermediate_17,
	intermediate_19,
	hps_io_usb1_inst_STP,
	intermediate_20,
	intermediate_22,
	intermediate_24,
	intermediate_26,
	intermediate_28,
	intermediate_30,
	intermediate_32,
	intermediate_34,
	intermediate_21,
	intermediate_23,
	intermediate_25,
	intermediate_27,
	intermediate_29,
	intermediate_31,
	intermediate_33,
	intermediate_35,
	hps_io_spim1_inst_CLK,
	hps_io_spim1_inst_SS0,
	intermediate_36,
	intermediate_37,
	hps_io_uart0_inst_TX,
	intermediate_39,
	intermediate_38,
	intermediate_41,
	intermediate_40,
	intermediate_42,
	intermediate_43,
	intermediate_44,
	intermediate_46,
	intermediate_48,
	intermediate_50,
	intermediate_52,
	intermediate_54,
	intermediate_45,
	intermediate_47,
	intermediate_49,
	intermediate_51,
	intermediate_53,
	intermediate_55,
	intermediate_56,
	intermediate_57,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_qspi_inst_IO0_0,
	hps_io_qspi_inst_IO1_0,
	hps_io_qspi_inst_IO2_0,
	hps_io_qspi_inst_IO3_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_io_usb1_inst_D0_0,
	hps_io_usb1_inst_D1_0,
	hps_io_usb1_inst_D2_0,
	hps_io_usb1_inst_D3_0,
	hps_io_usb1_inst_D4_0,
	hps_io_usb1_inst_D5_0,
	hps_io_usb1_inst_D6_0,
	hps_io_usb1_inst_D7_0,
	hps_io_i2c0_inst_SDA_0,
	hps_io_i2c0_inst_SCL_0,
	hps_io_i2c1_inst_SDA_0,
	hps_io_i2c1_inst_SCL_0,
	hps_io_gpio_inst_GPIO09_0,
	hps_io_gpio_inst_GPIO35_0,
	hps_io_gpio_inst_GPIO40_0,
	hps_io_gpio_inst_GPIO41_0,
	hps_io_gpio_inst_GPIO48_0,
	hps_io_gpio_inst_GPIO53_0,
	hps_io_gpio_inst_GPIO54_0,
	hps_io_gpio_inst_GPIO61_0,
	hps_io_emac1_inst_RXD0,
	hps_io_emac1_inst_RXD1,
	hps_io_emac1_inst_RXD2,
	hps_io_emac1_inst_RXD3,
	hps_io_emac1_inst_RX_CLK,
	hps_io_emac1_inst_RX_CTL,
	hps_io_spim1_inst_MISO,
	hps_io_uart0_inst_RX,
	hps_io_usb1_inst_CLK,
	hps_io_usb1_inst_DIR,
	hps_io_usb1_inst_NXT,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	[0:0] hps_io_emac1_inst_TX_CLK;
output 	[0:0] hps_io_emac1_inst_TX_CTL;
output 	intermediate_0;
output 	intermediate_1;
output 	[0:0] hps_io_emac1_inst_MDC;
output 	[0:0] hps_io_emac1_inst_TXD0;
output 	[0:0] hps_io_emac1_inst_TXD1;
output 	[0:0] hps_io_emac1_inst_TXD2;
output 	[0:0] hps_io_emac1_inst_TXD3;
output 	[0:0] hps_io_qspi_inst_CLK;
output 	intermediate_2;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_3;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	[0:0] hps_io_qspi_inst_SS0;
output 	[0:0] hps_io_sdio_inst_CLK;
output 	intermediate_10;
output 	intermediate_11;
output 	intermediate_12;
output 	intermediate_14;
output 	intermediate_16;
output 	intermediate_18;
output 	intermediate_13;
output 	intermediate_15;
output 	intermediate_17;
output 	intermediate_19;
output 	[0:0] hps_io_usb1_inst_STP;
output 	intermediate_20;
output 	intermediate_22;
output 	intermediate_24;
output 	intermediate_26;
output 	intermediate_28;
output 	intermediate_30;
output 	intermediate_32;
output 	intermediate_34;
output 	intermediate_21;
output 	intermediate_23;
output 	intermediate_25;
output 	intermediate_27;
output 	intermediate_29;
output 	intermediate_31;
output 	intermediate_33;
output 	intermediate_35;
output 	[0:0] hps_io_spim1_inst_CLK;
output 	[0:0] hps_io_spim1_inst_SS0;
output 	intermediate_36;
output 	intermediate_37;
output 	[0:0] hps_io_uart0_inst_TX;
output 	intermediate_39;
output 	intermediate_38;
output 	intermediate_41;
output 	intermediate_40;
output 	intermediate_42;
output 	intermediate_43;
output 	intermediate_44;
output 	intermediate_46;
output 	intermediate_48;
output 	intermediate_50;
output 	intermediate_52;
output 	intermediate_54;
output 	intermediate_45;
output 	intermediate_47;
output 	intermediate_49;
output 	intermediate_51;
output 	intermediate_53;
output 	intermediate_55;
output 	intermediate_56;
output 	intermediate_57;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_qspi_inst_IO0_0;
input 	hps_io_qspi_inst_IO1_0;
input 	hps_io_qspi_inst_IO2_0;
input 	hps_io_qspi_inst_IO3_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_io_usb1_inst_D0_0;
input 	hps_io_usb1_inst_D1_0;
input 	hps_io_usb1_inst_D2_0;
input 	hps_io_usb1_inst_D3_0;
input 	hps_io_usb1_inst_D4_0;
input 	hps_io_usb1_inst_D5_0;
input 	hps_io_usb1_inst_D6_0;
input 	hps_io_usb1_inst_D7_0;
input 	hps_io_i2c0_inst_SDA_0;
input 	hps_io_i2c0_inst_SCL_0;
input 	hps_io_i2c1_inst_SDA_0;
input 	hps_io_i2c1_inst_SCL_0;
input 	hps_io_gpio_inst_GPIO09_0;
input 	hps_io_gpio_inst_GPIO35_0;
input 	hps_io_gpio_inst_GPIO40_0;
input 	hps_io_gpio_inst_GPIO41_0;
input 	hps_io_gpio_inst_GPIO48_0;
input 	hps_io_gpio_inst_GPIO53_0;
input 	hps_io_gpio_inst_GPIO54_0;
input 	hps_io_gpio_inst_GPIO61_0;
input 	[0:0] hps_io_emac1_inst_RXD0;
input 	[0:0] hps_io_emac1_inst_RXD1;
input 	[0:0] hps_io_emac1_inst_RXD2;
input 	[0:0] hps_io_emac1_inst_RXD3;
input 	[0:0] hps_io_emac1_inst_RX_CLK;
input 	[0:0] hps_io_emac1_inst_RX_CTL;
input 	[0:0] hps_io_spim1_inst_MISO;
input 	[0:0] hps_io_uart0_inst_RX;
input 	[0:0] hps_io_usb1_inst_CLK;
input 	[0:0] hps_io_usb1_inst_DIR;
input 	[0:0] hps_io_usb1_inst_NXT;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sdio_inst~O_SDMMC_PWR_EN ;
wire \uart0_inst~UARTRTSN ;
wire \gpio_inst~LOANIO0_I0 ;
wire \gpio_inst~LOANIO0_I1 ;
wire \gpio_inst~LOANIO0_I2 ;
wire \gpio_inst~LOANIO0_I3 ;
wire \gpio_inst~LOANIO0_I4 ;
wire \gpio_inst~LOANIO0_I5 ;
wire \gpio_inst~LOANIO0_I6 ;
wire \gpio_inst~LOANIO0_I7 ;
wire \gpio_inst~LOANIO0_I8 ;
wire \gpio_inst~LOANIO0_I9 ;
wire \gpio_inst~LOANIO0_I10 ;
wire \gpio_inst~LOANIO0_I11 ;
wire \gpio_inst~LOANIO0_I12 ;
wire \gpio_inst~LOANIO0_I13 ;
wire \gpio_inst~LOANIO0_I14 ;
wire \gpio_inst~LOANIO0_I15 ;
wire \gpio_inst~LOANIO0_I16 ;
wire \gpio_inst~LOANIO0_I17 ;
wire \gpio_inst~LOANIO0_I18 ;
wire \gpio_inst~LOANIO0_I19 ;
wire \gpio_inst~LOANIO0_I20 ;
wire \gpio_inst~LOANIO0_I21 ;
wire \gpio_inst~LOANIO0_I22 ;
wire \gpio_inst~LOANIO0_I23 ;
wire \gpio_inst~LOANIO0_I24 ;
wire \gpio_inst~LOANIO0_I25 ;
wire \gpio_inst~LOANIO0_I26 ;
wire \gpio_inst~LOANIO0_I27 ;
wire \gpio_inst~LOANIO0_I28 ;
wire \~GND~combout ;

wire [3:0] emac1_inst_EMAC_PHY_TXD_bus;
wire [3:0] qspi_inst_QSPI_SS_N_bus;
wire [3:0] qspi_inst_QSPI_MO_EN_N_bus;
wire [7:0] sdio_inst_SDMMC_DATA_OE_bus;
wire [7:0] sdio_inst_SDMMC_DATA_O_bus;
wire [7:0] usb1_inst_USB_ULPI_DATA_O_bus;
wire [7:0] usb1_inst_USB_ULPI_DATA_OE_bus;
wire [28:0] gpio_inst_GPIO1_PORTA_O_bus;
wire [28:0] gpio_inst_GPIO0_PORTA_OE_bus;
wire [12:0] gpio_inst_GPIO2_PORTA_O_bus;
wire [28:0] gpio_inst_GPIO0_PORTA_O_bus;
wire [12:0] gpio_inst_GPIO2_PORTA_OE_bus;
wire [28:0] gpio_inst_GPIO1_PORTA_OE_bus;
wire [28:0] gpio_inst_LOANIO0_I_bus;

assign hps_io_emac1_inst_TXD0[0] = emac1_inst_EMAC_PHY_TXD_bus[0];
assign hps_io_emac1_inst_TXD1[0] = emac1_inst_EMAC_PHY_TXD_bus[1];
assign hps_io_emac1_inst_TXD2[0] = emac1_inst_EMAC_PHY_TXD_bus[2];
assign hps_io_emac1_inst_TXD3[0] = emac1_inst_EMAC_PHY_TXD_bus[3];

assign hps_io_qspi_inst_SS0[0] = qspi_inst_QSPI_SS_N_bus[0];

assign intermediate_3 = qspi_inst_QSPI_MO_EN_N_bus[0];
assign intermediate_5 = qspi_inst_QSPI_MO_EN_N_bus[1];
assign intermediate_7 = qspi_inst_QSPI_MO_EN_N_bus[2];
assign intermediate_9 = qspi_inst_QSPI_MO_EN_N_bus[3];

assign intermediate_13 = sdio_inst_SDMMC_DATA_OE_bus[0];
assign intermediate_15 = sdio_inst_SDMMC_DATA_OE_bus[1];
assign intermediate_17 = sdio_inst_SDMMC_DATA_OE_bus[2];
assign intermediate_19 = sdio_inst_SDMMC_DATA_OE_bus[3];

assign intermediate_12 = sdio_inst_SDMMC_DATA_O_bus[0];
assign intermediate_14 = sdio_inst_SDMMC_DATA_O_bus[1];
assign intermediate_16 = sdio_inst_SDMMC_DATA_O_bus[2];
assign intermediate_18 = sdio_inst_SDMMC_DATA_O_bus[3];

assign intermediate_20 = usb1_inst_USB_ULPI_DATA_O_bus[0];
assign intermediate_22 = usb1_inst_USB_ULPI_DATA_O_bus[1];
assign intermediate_24 = usb1_inst_USB_ULPI_DATA_O_bus[2];
assign intermediate_26 = usb1_inst_USB_ULPI_DATA_O_bus[3];
assign intermediate_28 = usb1_inst_USB_ULPI_DATA_O_bus[4];
assign intermediate_30 = usb1_inst_USB_ULPI_DATA_O_bus[5];
assign intermediate_32 = usb1_inst_USB_ULPI_DATA_O_bus[6];
assign intermediate_34 = usb1_inst_USB_ULPI_DATA_O_bus[7];

assign intermediate_21 = usb1_inst_USB_ULPI_DATA_OE_bus[0];
assign intermediate_23 = usb1_inst_USB_ULPI_DATA_OE_bus[1];
assign intermediate_25 = usb1_inst_USB_ULPI_DATA_OE_bus[2];
assign intermediate_27 = usb1_inst_USB_ULPI_DATA_OE_bus[3];
assign intermediate_29 = usb1_inst_USB_ULPI_DATA_OE_bus[4];
assign intermediate_31 = usb1_inst_USB_ULPI_DATA_OE_bus[5];
assign intermediate_33 = usb1_inst_USB_ULPI_DATA_OE_bus[6];
assign intermediate_35 = usb1_inst_USB_ULPI_DATA_OE_bus[7];

assign intermediate_44 = gpio_inst_GPIO1_PORTA_O_bus[6];
assign intermediate_46 = gpio_inst_GPIO1_PORTA_O_bus[11];
assign intermediate_48 = gpio_inst_GPIO1_PORTA_O_bus[12];
assign intermediate_50 = gpio_inst_GPIO1_PORTA_O_bus[19];
assign intermediate_52 = gpio_inst_GPIO1_PORTA_O_bus[24];
assign intermediate_54 = gpio_inst_GPIO1_PORTA_O_bus[25];

assign intermediate_43 = gpio_inst_GPIO0_PORTA_OE_bus[9];

assign intermediate_56 = gpio_inst_GPIO2_PORTA_O_bus[3];

assign intermediate_42 = gpio_inst_GPIO0_PORTA_O_bus[9];

assign intermediate_57 = gpio_inst_GPIO2_PORTA_OE_bus[3];

assign intermediate_45 = gpio_inst_GPIO1_PORTA_OE_bus[6];
assign intermediate_47 = gpio_inst_GPIO1_PORTA_OE_bus[11];
assign intermediate_49 = gpio_inst_GPIO1_PORTA_OE_bus[12];
assign intermediate_51 = gpio_inst_GPIO1_PORTA_OE_bus[19];
assign intermediate_53 = gpio_inst_GPIO1_PORTA_OE_bus[24];
assign intermediate_55 = gpio_inst_GPIO1_PORTA_OE_bus[25];

assign \gpio_inst~LOANIO0_I0  = gpio_inst_LOANIO0_I_bus[0];
assign \gpio_inst~LOANIO0_I1  = gpio_inst_LOANIO0_I_bus[1];
assign \gpio_inst~LOANIO0_I2  = gpio_inst_LOANIO0_I_bus[2];
assign \gpio_inst~LOANIO0_I3  = gpio_inst_LOANIO0_I_bus[3];
assign \gpio_inst~LOANIO0_I4  = gpio_inst_LOANIO0_I_bus[4];
assign \gpio_inst~LOANIO0_I5  = gpio_inst_LOANIO0_I_bus[5];
assign \gpio_inst~LOANIO0_I6  = gpio_inst_LOANIO0_I_bus[6];
assign \gpio_inst~LOANIO0_I7  = gpio_inst_LOANIO0_I_bus[7];
assign \gpio_inst~LOANIO0_I8  = gpio_inst_LOANIO0_I_bus[8];
assign \gpio_inst~LOANIO0_I9  = gpio_inst_LOANIO0_I_bus[9];
assign \gpio_inst~LOANIO0_I10  = gpio_inst_LOANIO0_I_bus[10];
assign \gpio_inst~LOANIO0_I11  = gpio_inst_LOANIO0_I_bus[11];
assign \gpio_inst~LOANIO0_I12  = gpio_inst_LOANIO0_I_bus[12];
assign \gpio_inst~LOANIO0_I13  = gpio_inst_LOANIO0_I_bus[13];
assign \gpio_inst~LOANIO0_I14  = gpio_inst_LOANIO0_I_bus[14];
assign \gpio_inst~LOANIO0_I15  = gpio_inst_LOANIO0_I_bus[15];
assign \gpio_inst~LOANIO0_I16  = gpio_inst_LOANIO0_I_bus[16];
assign \gpio_inst~LOANIO0_I17  = gpio_inst_LOANIO0_I_bus[17];
assign \gpio_inst~LOANIO0_I18  = gpio_inst_LOANIO0_I_bus[18];
assign \gpio_inst~LOANIO0_I19  = gpio_inst_LOANIO0_I_bus[19];
assign \gpio_inst~LOANIO0_I20  = gpio_inst_LOANIO0_I_bus[20];
assign \gpio_inst~LOANIO0_I21  = gpio_inst_LOANIO0_I_bus[21];
assign \gpio_inst~LOANIO0_I22  = gpio_inst_LOANIO0_I_bus[22];
assign \gpio_inst~LOANIO0_I23  = gpio_inst_LOANIO0_I_bus[23];
assign \gpio_inst~LOANIO0_I24  = gpio_inst_LOANIO0_I_bus[24];
assign \gpio_inst~LOANIO0_I25  = gpio_inst_LOANIO0_I_bus[25];
assign \gpio_inst~LOANIO0_I26  = gpio_inst_LOANIO0_I_bus[26];
assign \gpio_inst~LOANIO0_I27  = gpio_inst_LOANIO0_I_bus[27];
assign \gpio_inst~LOANIO0_I28  = gpio_inst_LOANIO0_I_bus[28];

Computer_System_hps_sdram hps_sdram_inst(
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.GND_port(\~GND~combout ),
	.memory_oct_rzqin(memory_oct_rzqin));

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

cyclonev_hps_peripheral_emac emac1_inst(
	.emac_clk_rx(hps_io_emac1_inst_RX_CLK[0]),
	.emac_phy_rxdv(hps_io_emac1_inst_RX_CTL[0]),
	.emac_gmii_mdo_i(hps_io_emac1_inst_MDIO_0),
	.emac_phy_rxd({hps_io_emac1_inst_RXD3[0],hps_io_emac1_inst_RXD2[0],hps_io_emac1_inst_RXD1[0],hps_io_emac1_inst_RXD0[0]}),
	.emac_clk_tx(hps_io_emac1_inst_TX_CLK[0]),
	.emac_phy_tx_oe(hps_io_emac1_inst_TX_CTL[0]),
	.emac_gmii_mdo_o(intermediate_0),
	.emac_gmii_mdo_oe(intermediate_1),
	.emac_gmii_mdc(hps_io_emac1_inst_MDC[0]),
	.emac_phy_txd(emac1_inst_EMAC_PHY_TXD_bus));
defparam emac1_inst.dummy_param = 256;

cyclonev_hps_peripheral_qspi qspi_inst(
	.qspi_mi0(hps_io_qspi_inst_IO0_0),
	.qspi_mi1(hps_io_qspi_inst_IO1_0),
	.qspi_mi2(hps_io_qspi_inst_IO2_0),
	.qspi_mi3(hps_io_qspi_inst_IO3_0),
	.qspi_sclk(hps_io_qspi_inst_CLK[0]),
	.qspi_mo0(intermediate_2),
	.qspi_mo1(intermediate_4),
	.qspi_mo2(intermediate_6),
	.qspi_mo3(intermediate_8),
	.qspi_mo_en_n(qspi_inst_QSPI_MO_EN_N_bus),
	.qspi_ss_n(qspi_inst_QSPI_SS_N_bus));
defparam qspi_inst.dummy_param = 256;

cyclonev_hps_peripheral_sdmmc sdio_inst(
	.sdmmc_fb_clk(gnd),
	.sdmmc_cmd_i(hps_io_sdio_inst_CMD_0),
	.sdmmc_data_i({gnd,gnd,gnd,gnd,hps_io_sdio_inst_D3_0,hps_io_sdio_inst_D2_0,hps_io_sdio_inst_D1_0,hps_io_sdio_inst_D0_0}),
	.sdmmc_pwr_en(\sdio_inst~O_SDMMC_PWR_EN ),
	.sdmmc_cclk(hps_io_sdio_inst_CLK[0]),
	.sdmmc_cmd_o(intermediate_10),
	.sdmmc_cmd_oe(intermediate_11),
	.sdmmc_data_o(sdio_inst_SDMMC_DATA_O_bus),
	.sdmmc_data_oe(sdio_inst_SDMMC_DATA_OE_bus));
defparam sdio_inst.dummy_param = 256;

cyclonev_hps_peripheral_usb usb1_inst(
	.usb_ulpi_clk(hps_io_usb1_inst_CLK[0]),
	.usb_ulpi_dir(hps_io_usb1_inst_DIR[0]),
	.usb_ulpi_nxt(hps_io_usb1_inst_NXT[0]),
	.usb_ulpi_data_i({hps_io_usb1_inst_D7_0,hps_io_usb1_inst_D6_0,hps_io_usb1_inst_D5_0,hps_io_usb1_inst_D4_0,hps_io_usb1_inst_D3_0,hps_io_usb1_inst_D2_0,hps_io_usb1_inst_D1_0,hps_io_usb1_inst_D0_0}),
	.usb_ulpi_stp(hps_io_usb1_inst_STP[0]),
	.usb_ulpi_data_o(usb1_inst_USB_ULPI_DATA_O_bus),
	.usb_ulpi_data_oe(usb1_inst_USB_ULPI_DATA_OE_bus));
defparam usb1_inst.dummy_param = 256;

cyclonev_hps_peripheral_spi_master spim1_inst(
	.spi_master_rxd(hps_io_spim1_inst_MISO[0]),
	.spi_master_sclk(hps_io_spim1_inst_CLK[0]),
	.spi_master_ss_0_n(hps_io_spim1_inst_SS0[0]),
	.spi_master_ss_1_n(),
	.spi_master_txd(intermediate_36),
	.spi_master_ssi_oe_n(intermediate_37));
defparam spim1_inst.dummy_param = 256;

cyclonev_hps_peripheral_uart uart0_inst(
	.uart_cts_n(gnd),
	.uart_rxd(hps_io_uart0_inst_RX[0]),
	.uart_rts_n(\uart0_inst~UARTRTSN ),
	.uart_txd(hps_io_uart0_inst_TX[0]));
defparam uart0_inst.dummy_param = 256;

cyclonev_hps_peripheral_i2c i2c0_inst(
	.i2c_clk(hps_io_i2c0_inst_SCL_0),
	.i2c_data(hps_io_i2c0_inst_SDA_0),
	.i2c_clk_oe(intermediate_39),
	.i2c_data_oe(intermediate_38));
defparam i2c0_inst.dummy_param = 256;

cyclonev_hps_peripheral_i2c i2c1_inst(
	.i2c_clk(hps_io_i2c1_inst_SCL_0),
	.i2c_data(hps_io_i2c1_inst_SDA_0),
	.i2c_clk_oe(intermediate_41),
	.i2c_data_oe(intermediate_40));
defparam i2c1_inst.dummy_param = 256;

cyclonev_hps_peripheral_gpio gpio_inst(
	.gpio0_porta_i({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,hps_io_gpio_inst_GPIO09_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.gpio1_porta_i({gnd,gnd,gnd,hps_io_gpio_inst_GPIO54_0,hps_io_gpio_inst_GPIO53_0,gnd,gnd,gnd,gnd,hps_io_gpio_inst_GPIO48_0,gnd,gnd,gnd,gnd,gnd,gnd,hps_io_gpio_inst_GPIO41_0,hps_io_gpio_inst_GPIO40_0,gnd,gnd,gnd,gnd,hps_io_gpio_inst_GPIO35_0,gnd,gnd,gnd,gnd,gnd,gnd}),
	.gpio2_porta_i({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,hps_io_gpio_inst_GPIO61_0,gnd,gnd,gnd}),
	.loanio0_o(29'b00000000000000000000000000000),
	.loanio0_oe(29'b00000000000000000000000000000),
	.loanio1_o(29'b00000000000000000000000000000),
	.loanio1_oe(29'b00000000000000000000000000000),
	.loanio2_o(29'b00000000000000000000000000000),
	.loanio2_oe(29'b00000000000000000000000000000),
	.loanio0_i(gpio_inst_LOANIO0_I_bus),
	.loanio1_i(),
	.loanio2_i(),
	.gpio0_porta_o(gpio_inst_GPIO0_PORTA_O_bus),
	.gpio0_porta_oe(gpio_inst_GPIO0_PORTA_OE_bus),
	.gpio1_porta_o(gpio_inst_GPIO1_PORTA_O_bus),
	.gpio1_porta_oe(gpio_inst_GPIO1_PORTA_OE_bus),
	.gpio2_porta_o(gpio_inst_GPIO2_PORTA_O_bus),
	.gpio2_porta_oe(gpio_inst_GPIO2_PORTA_OE_bus));
defparam gpio_inst.dummy_param = 256;

endmodule

module Computer_System_hps_sdram (
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	GND_port,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	GND_port;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \pll|afi_clk ;
wire \pll|pll_write_clk ;
wire \p0|umemphy|afi_cal_fail ;
wire \p0|umemphy|afi_cal_success ;
wire \p0|umemphy|afi_rdata_valid[0] ;
wire \p0|umemphy|ctl_reset_n ;
wire \p0|umemphy|afi_rdata[0] ;
wire \p0|umemphy|afi_rdata[1] ;
wire \p0|umemphy|afi_rdata[2] ;
wire \p0|umemphy|afi_rdata[3] ;
wire \p0|umemphy|afi_rdata[4] ;
wire \p0|umemphy|afi_rdata[5] ;
wire \p0|umemphy|afi_rdata[6] ;
wire \p0|umemphy|afi_rdata[7] ;
wire \p0|umemphy|afi_rdata[8] ;
wire \p0|umemphy|afi_rdata[9] ;
wire \p0|umemphy|afi_rdata[10] ;
wire \p0|umemphy|afi_rdata[11] ;
wire \p0|umemphy|afi_rdata[12] ;
wire \p0|umemphy|afi_rdata[13] ;
wire \p0|umemphy|afi_rdata[14] ;
wire \p0|umemphy|afi_rdata[15] ;
wire \p0|umemphy|afi_rdata[16] ;
wire \p0|umemphy|afi_rdata[17] ;
wire \p0|umemphy|afi_rdata[18] ;
wire \p0|umemphy|afi_rdata[19] ;
wire \p0|umemphy|afi_rdata[20] ;
wire \p0|umemphy|afi_rdata[21] ;
wire \p0|umemphy|afi_rdata[22] ;
wire \p0|umemphy|afi_rdata[23] ;
wire \p0|umemphy|afi_rdata[24] ;
wire \p0|umemphy|afi_rdata[25] ;
wire \p0|umemphy|afi_rdata[26] ;
wire \p0|umemphy|afi_rdata[27] ;
wire \p0|umemphy|afi_rdata[28] ;
wire \p0|umemphy|afi_rdata[29] ;
wire \p0|umemphy|afi_rdata[30] ;
wire \p0|umemphy|afi_rdata[31] ;
wire \p0|umemphy|afi_rdata[32] ;
wire \p0|umemphy|afi_rdata[33] ;
wire \p0|umemphy|afi_rdata[34] ;
wire \p0|umemphy|afi_rdata[35] ;
wire \p0|umemphy|afi_rdata[36] ;
wire \p0|umemphy|afi_rdata[37] ;
wire \p0|umemphy|afi_rdata[38] ;
wire \p0|umemphy|afi_rdata[39] ;
wire \p0|umemphy|afi_rdata[40] ;
wire \p0|umemphy|afi_rdata[41] ;
wire \p0|umemphy|afi_rdata[42] ;
wire \p0|umemphy|afi_rdata[43] ;
wire \p0|umemphy|afi_rdata[44] ;
wire \p0|umemphy|afi_rdata[45] ;
wire \p0|umemphy|afi_rdata[46] ;
wire \p0|umemphy|afi_rdata[47] ;
wire \p0|umemphy|afi_rdata[48] ;
wire \p0|umemphy|afi_rdata[49] ;
wire \p0|umemphy|afi_rdata[50] ;
wire \p0|umemphy|afi_rdata[51] ;
wire \p0|umemphy|afi_rdata[52] ;
wire \p0|umemphy|afi_rdata[53] ;
wire \p0|umemphy|afi_rdata[54] ;
wire \p0|umemphy|afi_rdata[55] ;
wire \p0|umemphy|afi_rdata[56] ;
wire \p0|umemphy|afi_rdata[57] ;
wire \p0|umemphy|afi_rdata[58] ;
wire \p0|umemphy|afi_rdata[59] ;
wire \p0|umemphy|afi_rdata[60] ;
wire \p0|umemphy|afi_rdata[61] ;
wire \p0|umemphy|afi_rdata[62] ;
wire \p0|umemphy|afi_rdata[63] ;
wire \p0|umemphy|afi_rdata[64] ;
wire \p0|umemphy|afi_rdata[65] ;
wire \p0|umemphy|afi_rdata[66] ;
wire \p0|umemphy|afi_rdata[67] ;
wire \p0|umemphy|afi_rdata[68] ;
wire \p0|umemphy|afi_rdata[69] ;
wire \p0|umemphy|afi_rdata[70] ;
wire \p0|umemphy|afi_rdata[71] ;
wire \p0|umemphy|afi_rdata[72] ;
wire \p0|umemphy|afi_rdata[73] ;
wire \p0|umemphy|afi_rdata[74] ;
wire \p0|umemphy|afi_rdata[75] ;
wire \p0|umemphy|afi_rdata[76] ;
wire \p0|umemphy|afi_rdata[77] ;
wire \p0|umemphy|afi_rdata[78] ;
wire \p0|umemphy|afi_rdata[79] ;
wire \p0|umemphy|afi_wlat[0] ;
wire \p0|umemphy|afi_wlat[1] ;
wire \p0|umemphy|afi_wlat[2] ;
wire \p0|umemphy|afi_wlat[3] ;
wire \c0|afi_cas_n[0] ;
wire \c0|afi_ras_n[0] ;
wire \c0|afi_rst_n[0] ;
wire \c0|afi_we_n[0] ;
wire \c0|afi_addr[0] ;
wire \c0|afi_addr[1] ;
wire \c0|afi_addr[2] ;
wire \c0|afi_addr[3] ;
wire \c0|afi_addr[4] ;
wire \c0|afi_addr[5] ;
wire \c0|afi_addr[6] ;
wire \c0|afi_addr[7] ;
wire \c0|afi_addr[8] ;
wire \c0|afi_addr[9] ;
wire \c0|afi_addr[10] ;
wire \c0|afi_addr[11] ;
wire \c0|afi_addr[12] ;
wire \c0|afi_addr[13] ;
wire \c0|afi_addr[14] ;
wire \c0|afi_addr[15] ;
wire \c0|afi_addr[16] ;
wire \c0|afi_addr[17] ;
wire \c0|afi_addr[18] ;
wire \c0|afi_addr[19] ;
wire \c0|afi_ba[0] ;
wire \c0|afi_ba[1] ;
wire \c0|afi_ba[2] ;
wire \c0|afi_cke[0] ;
wire \c0|afi_cke[1] ;
wire \c0|afi_cs_n[0] ;
wire \c0|afi_cs_n[1] ;
wire \c0|afi_dm_int[0] ;
wire \c0|afi_dm_int[1] ;
wire \c0|afi_dm_int[2] ;
wire \c0|afi_dm_int[3] ;
wire \c0|afi_dm_int[4] ;
wire \c0|afi_dm_int[5] ;
wire \c0|afi_dm_int[6] ;
wire \c0|afi_dm_int[7] ;
wire \c0|afi_dm_int[8] ;
wire \c0|afi_dm_int[9] ;
wire \c0|afi_dqs_burst[0] ;
wire \c0|afi_dqs_burst[1] ;
wire \c0|afi_dqs_burst[2] ;
wire \c0|afi_dqs_burst[3] ;
wire \c0|afi_dqs_burst[4] ;
wire \c0|afi_odt[0] ;
wire \c0|afi_odt[1] ;
wire \c0|afi_rdata_en[0] ;
wire \c0|afi_rdata_en[1] ;
wire \c0|afi_rdata_en[2] ;
wire \c0|afi_rdata_en[3] ;
wire \c0|afi_rdata_en[4] ;
wire \c0|afi_rdata_en_full[0] ;
wire \c0|afi_rdata_en_full[1] ;
wire \c0|afi_rdata_en_full[2] ;
wire \c0|afi_rdata_en_full[3] ;
wire \c0|afi_rdata_en_full[4] ;
wire \c0|afi_wdata_int[0] ;
wire \c0|afi_wdata_int[1] ;
wire \c0|afi_wdata_int[2] ;
wire \c0|afi_wdata_int[3] ;
wire \c0|afi_wdata_int[4] ;
wire \c0|afi_wdata_int[5] ;
wire \c0|afi_wdata_int[6] ;
wire \c0|afi_wdata_int[7] ;
wire \c0|afi_wdata_int[8] ;
wire \c0|afi_wdata_int[9] ;
wire \c0|afi_wdata_int[10] ;
wire \c0|afi_wdata_int[11] ;
wire \c0|afi_wdata_int[12] ;
wire \c0|afi_wdata_int[13] ;
wire \c0|afi_wdata_int[14] ;
wire \c0|afi_wdata_int[15] ;
wire \c0|afi_wdata_int[16] ;
wire \c0|afi_wdata_int[17] ;
wire \c0|afi_wdata_int[18] ;
wire \c0|afi_wdata_int[19] ;
wire \c0|afi_wdata_int[20] ;
wire \c0|afi_wdata_int[21] ;
wire \c0|afi_wdata_int[22] ;
wire \c0|afi_wdata_int[23] ;
wire \c0|afi_wdata_int[24] ;
wire \c0|afi_wdata_int[25] ;
wire \c0|afi_wdata_int[26] ;
wire \c0|afi_wdata_int[27] ;
wire \c0|afi_wdata_int[28] ;
wire \c0|afi_wdata_int[29] ;
wire \c0|afi_wdata_int[30] ;
wire \c0|afi_wdata_int[31] ;
wire \c0|afi_wdata_int[32] ;
wire \c0|afi_wdata_int[33] ;
wire \c0|afi_wdata_int[34] ;
wire \c0|afi_wdata_int[35] ;
wire \c0|afi_wdata_int[36] ;
wire \c0|afi_wdata_int[37] ;
wire \c0|afi_wdata_int[38] ;
wire \c0|afi_wdata_int[39] ;
wire \c0|afi_wdata_int[40] ;
wire \c0|afi_wdata_int[41] ;
wire \c0|afi_wdata_int[42] ;
wire \c0|afi_wdata_int[43] ;
wire \c0|afi_wdata_int[44] ;
wire \c0|afi_wdata_int[45] ;
wire \c0|afi_wdata_int[46] ;
wire \c0|afi_wdata_int[47] ;
wire \c0|afi_wdata_int[48] ;
wire \c0|afi_wdata_int[49] ;
wire \c0|afi_wdata_int[50] ;
wire \c0|afi_wdata_int[51] ;
wire \c0|afi_wdata_int[52] ;
wire \c0|afi_wdata_int[53] ;
wire \c0|afi_wdata_int[54] ;
wire \c0|afi_wdata_int[55] ;
wire \c0|afi_wdata_int[56] ;
wire \c0|afi_wdata_int[57] ;
wire \c0|afi_wdata_int[58] ;
wire \c0|afi_wdata_int[59] ;
wire \c0|afi_wdata_int[60] ;
wire \c0|afi_wdata_int[61] ;
wire \c0|afi_wdata_int[62] ;
wire \c0|afi_wdata_int[63] ;
wire \c0|afi_wdata_int[64] ;
wire \c0|afi_wdata_int[65] ;
wire \c0|afi_wdata_int[66] ;
wire \c0|afi_wdata_int[67] ;
wire \c0|afi_wdata_int[68] ;
wire \c0|afi_wdata_int[69] ;
wire \c0|afi_wdata_int[70] ;
wire \c0|afi_wdata_int[71] ;
wire \c0|afi_wdata_int[72] ;
wire \c0|afi_wdata_int[73] ;
wire \c0|afi_wdata_int[74] ;
wire \c0|afi_wdata_int[75] ;
wire \c0|afi_wdata_int[76] ;
wire \c0|afi_wdata_int[77] ;
wire \c0|afi_wdata_int[78] ;
wire \c0|afi_wdata_int[79] ;
wire \c0|afi_wdata_valid[0] ;
wire \c0|afi_wdata_valid[1] ;
wire \c0|afi_wdata_valid[2] ;
wire \c0|afi_wdata_valid[3] ;
wire \c0|afi_wdata_valid[4] ;
wire \c0|cfg_addlat_wire[0] ;
wire \c0|cfg_addlat_wire[1] ;
wire \c0|cfg_addlat_wire[2] ;
wire \c0|cfg_addlat_wire[3] ;
wire \c0|cfg_addlat_wire[4] ;
wire \c0|cfg_bankaddrwidth_wire[0] ;
wire \c0|cfg_bankaddrwidth_wire[1] ;
wire \c0|cfg_bankaddrwidth_wire[2] ;
wire \c0|cfg_caswrlat_wire[0] ;
wire \c0|cfg_caswrlat_wire[1] ;
wire \c0|cfg_caswrlat_wire[2] ;
wire \c0|cfg_caswrlat_wire[3] ;
wire \c0|cfg_coladdrwidth_wire[0] ;
wire \c0|cfg_coladdrwidth_wire[1] ;
wire \c0|cfg_coladdrwidth_wire[2] ;
wire \c0|cfg_coladdrwidth_wire[3] ;
wire \c0|cfg_coladdrwidth_wire[4] ;
wire \c0|cfg_csaddrwidth_wire[0] ;
wire \c0|cfg_csaddrwidth_wire[1] ;
wire \c0|cfg_csaddrwidth_wire[2] ;
wire \c0|cfg_devicewidth_wire[0] ;
wire \c0|cfg_devicewidth_wire[1] ;
wire \c0|cfg_devicewidth_wire[2] ;
wire \c0|cfg_devicewidth_wire[3] ;
wire \c0|cfg_interfacewidth_wire[0] ;
wire \c0|cfg_interfacewidth_wire[1] ;
wire \c0|cfg_interfacewidth_wire[2] ;
wire \c0|cfg_interfacewidth_wire[3] ;
wire \c0|cfg_interfacewidth_wire[4] ;
wire \c0|cfg_interfacewidth_wire[5] ;
wire \c0|cfg_interfacewidth_wire[6] ;
wire \c0|cfg_interfacewidth_wire[7] ;
wire \c0|cfg_rowaddrwidth_wire[0] ;
wire \c0|cfg_rowaddrwidth_wire[1] ;
wire \c0|cfg_rowaddrwidth_wire[2] ;
wire \c0|cfg_rowaddrwidth_wire[3] ;
wire \c0|cfg_rowaddrwidth_wire[4] ;
wire \c0|cfg_tcl_wire[0] ;
wire \c0|cfg_tcl_wire[1] ;
wire \c0|cfg_tcl_wire[2] ;
wire \c0|cfg_tcl_wire[3] ;
wire \c0|cfg_tcl_wire[4] ;
wire \c0|cfg_tmrd_wire[0] ;
wire \c0|cfg_tmrd_wire[1] ;
wire \c0|cfg_tmrd_wire[2] ;
wire \c0|cfg_tmrd_wire[3] ;
wire \c0|cfg_trefi_wire[0] ;
wire \c0|cfg_trefi_wire[1] ;
wire \c0|cfg_trefi_wire[2] ;
wire \c0|cfg_trefi_wire[3] ;
wire \c0|cfg_trefi_wire[4] ;
wire \c0|cfg_trefi_wire[5] ;
wire \c0|cfg_trefi_wire[6] ;
wire \c0|cfg_trefi_wire[7] ;
wire \c0|cfg_trefi_wire[8] ;
wire \c0|cfg_trefi_wire[9] ;
wire \c0|cfg_trefi_wire[10] ;
wire \c0|cfg_trefi_wire[11] ;
wire \c0|cfg_trefi_wire[12] ;
wire \c0|cfg_trfc_wire[0] ;
wire \c0|cfg_trfc_wire[1] ;
wire \c0|cfg_trfc_wire[2] ;
wire \c0|cfg_trfc_wire[3] ;
wire \c0|cfg_trfc_wire[4] ;
wire \c0|cfg_trfc_wire[5] ;
wire \c0|cfg_trfc_wire[6] ;
wire \c0|cfg_trfc_wire[7] ;
wire \c0|cfg_twr_wire[0] ;
wire \c0|cfg_twr_wire[1] ;
wire \c0|cfg_twr_wire[2] ;
wire \c0|cfg_twr_wire[3] ;
wire \c0|afi_mem_clk_disable[0] ;
wire \c0|cfg_dramconfig_wire[0] ;
wire \c0|cfg_dramconfig_wire[1] ;
wire \c0|cfg_dramconfig_wire[2] ;
wire \c0|cfg_dramconfig_wire[3] ;
wire \c0|cfg_dramconfig_wire[4] ;
wire \c0|cfg_dramconfig_wire[5] ;
wire \c0|cfg_dramconfig_wire[6] ;
wire \c0|cfg_dramconfig_wire[7] ;
wire \c0|cfg_dramconfig_wire[8] ;
wire \c0|cfg_dramconfig_wire[9] ;
wire \c0|cfg_dramconfig_wire[10] ;
wire \c0|cfg_dramconfig_wire[11] ;
wire \c0|cfg_dramconfig_wire[12] ;
wire \c0|cfg_dramconfig_wire[13] ;
wire \c0|cfg_dramconfig_wire[14] ;
wire \c0|cfg_dramconfig_wire[15] ;
wire \c0|cfg_dramconfig_wire[16] ;
wire \c0|cfg_dramconfig_wire[17] ;
wire \c0|cfg_dramconfig_wire[18] ;
wire \c0|cfg_dramconfig_wire[19] ;
wire \c0|cfg_dramconfig_wire[20] ;
wire \p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ;
wire \dll|dll_delayctrl[0] ;
wire \dll|dll_delayctrl[1] ;
wire \dll|dll_delayctrl[2] ;
wire \dll|dll_delayctrl[3] ;
wire \dll|dll_delayctrl[4] ;
wire \dll|dll_delayctrl[5] ;
wire \dll|dll_delayctrl[6] ;


Computer_System_altera_mem_if_dll_cyclonev dll(
	.clk(\pll|pll_write_clk ),
	.dll_delayctrl({\dll|dll_delayctrl[6] ,\dll|dll_delayctrl[5] ,\dll|dll_delayctrl[4] ,\dll|dll_delayctrl[3] ,\dll|dll_delayctrl[2] ,\dll|dll_delayctrl[1] ,\dll|dll_delayctrl[0] }));

Computer_System_altera_mem_if_oct_cyclonev oct(
	.parallelterminationcontrol({parallelterminationcontrol_15,parallelterminationcontrol_14,parallelterminationcontrol_13,parallelterminationcontrol_12,parallelterminationcontrol_11,parallelterminationcontrol_10,parallelterminationcontrol_9,parallelterminationcontrol_8,
parallelterminationcontrol_7,parallelterminationcontrol_6,parallelterminationcontrol_5,parallelterminationcontrol_4,parallelterminationcontrol_3,parallelterminationcontrol_2,parallelterminationcontrol_1,parallelterminationcontrol_0}),
	.seriesterminationcontrol({seriesterminationcontrol_15,seriesterminationcontrol_14,seriesterminationcontrol_13,seriesterminationcontrol_12,seriesterminationcontrol_11,seriesterminationcontrol_10,seriesterminationcontrol_9,seriesterminationcontrol_8,seriesterminationcontrol_7,
seriesterminationcontrol_6,seriesterminationcontrol_5,seriesterminationcontrol_4,seriesterminationcontrol_3,seriesterminationcontrol_2,seriesterminationcontrol_1,seriesterminationcontrol_0}),
	.oct_rzqin(memory_oct_rzqin));

Computer_System_altera_mem_if_hard_memory_controller_top_cyclonev c0(
	.afi_cal_fail(\p0|umemphy|afi_cal_fail ),
	.afi_cal_success(\p0|umemphy|afi_cal_success ),
	.afi_rdata_valid({\p0|umemphy|afi_rdata_valid[0] }),
	.ctl_reset_n(\p0|umemphy|ctl_reset_n ),
	.afi_rdata({\p0|umemphy|afi_rdata[79] ,\p0|umemphy|afi_rdata[78] ,\p0|umemphy|afi_rdata[77] ,\p0|umemphy|afi_rdata[76] ,\p0|umemphy|afi_rdata[75] ,\p0|umemphy|afi_rdata[74] ,\p0|umemphy|afi_rdata[73] ,\p0|umemphy|afi_rdata[72] ,\p0|umemphy|afi_rdata[71] ,
\p0|umemphy|afi_rdata[70] ,\p0|umemphy|afi_rdata[69] ,\p0|umemphy|afi_rdata[68] ,\p0|umemphy|afi_rdata[67] ,\p0|umemphy|afi_rdata[66] ,\p0|umemphy|afi_rdata[65] ,\p0|umemphy|afi_rdata[64] ,\p0|umemphy|afi_rdata[63] ,\p0|umemphy|afi_rdata[62] ,
\p0|umemphy|afi_rdata[61] ,\p0|umemphy|afi_rdata[60] ,\p0|umemphy|afi_rdata[59] ,\p0|umemphy|afi_rdata[58] ,\p0|umemphy|afi_rdata[57] ,\p0|umemphy|afi_rdata[56] ,\p0|umemphy|afi_rdata[55] ,\p0|umemphy|afi_rdata[54] ,\p0|umemphy|afi_rdata[53] ,
\p0|umemphy|afi_rdata[52] ,\p0|umemphy|afi_rdata[51] ,\p0|umemphy|afi_rdata[50] ,\p0|umemphy|afi_rdata[49] ,\p0|umemphy|afi_rdata[48] ,\p0|umemphy|afi_rdata[47] ,\p0|umemphy|afi_rdata[46] ,\p0|umemphy|afi_rdata[45] ,\p0|umemphy|afi_rdata[44] ,
\p0|umemphy|afi_rdata[43] ,\p0|umemphy|afi_rdata[42] ,\p0|umemphy|afi_rdata[41] ,\p0|umemphy|afi_rdata[40] ,\p0|umemphy|afi_rdata[39] ,\p0|umemphy|afi_rdata[38] ,\p0|umemphy|afi_rdata[37] ,\p0|umemphy|afi_rdata[36] ,\p0|umemphy|afi_rdata[35] ,
\p0|umemphy|afi_rdata[34] ,\p0|umemphy|afi_rdata[33] ,\p0|umemphy|afi_rdata[32] ,\p0|umemphy|afi_rdata[31] ,\p0|umemphy|afi_rdata[30] ,\p0|umemphy|afi_rdata[29] ,\p0|umemphy|afi_rdata[28] ,\p0|umemphy|afi_rdata[27] ,\p0|umemphy|afi_rdata[26] ,
\p0|umemphy|afi_rdata[25] ,\p0|umemphy|afi_rdata[24] ,\p0|umemphy|afi_rdata[23] ,\p0|umemphy|afi_rdata[22] ,\p0|umemphy|afi_rdata[21] ,\p0|umemphy|afi_rdata[20] ,\p0|umemphy|afi_rdata[19] ,\p0|umemphy|afi_rdata[18] ,\p0|umemphy|afi_rdata[17] ,
\p0|umemphy|afi_rdata[16] ,\p0|umemphy|afi_rdata[15] ,\p0|umemphy|afi_rdata[14] ,\p0|umemphy|afi_rdata[13] ,\p0|umemphy|afi_rdata[12] ,\p0|umemphy|afi_rdata[11] ,\p0|umemphy|afi_rdata[10] ,\p0|umemphy|afi_rdata[9] ,\p0|umemphy|afi_rdata[8] ,
\p0|umemphy|afi_rdata[7] ,\p0|umemphy|afi_rdata[6] ,\p0|umemphy|afi_rdata[5] ,\p0|umemphy|afi_rdata[4] ,\p0|umemphy|afi_rdata[3] ,\p0|umemphy|afi_rdata[2] ,\p0|umemphy|afi_rdata[1] ,\p0|umemphy|afi_rdata[0] }),
	.afi_wlat({\p0|umemphy|afi_wlat[3] ,\p0|umemphy|afi_wlat[2] ,\p0|umemphy|afi_wlat[1] ,\p0|umemphy|afi_wlat[0] }),
	.afi_cas_n({\c0|afi_cas_n[0] }),
	.afi_ras_n({\c0|afi_ras_n[0] }),
	.afi_rst_n({\c0|afi_rst_n[0] }),
	.afi_we_n({\c0|afi_we_n[0] }),
	.afi_addr({\c0|afi_addr[19] ,\c0|afi_addr[18] ,\c0|afi_addr[17] ,\c0|afi_addr[16] ,\c0|afi_addr[15] ,\c0|afi_addr[14] ,\c0|afi_addr[13] ,\c0|afi_addr[12] ,\c0|afi_addr[11] ,\c0|afi_addr[10] ,\c0|afi_addr[9] ,\c0|afi_addr[8] ,\c0|afi_addr[7] ,\c0|afi_addr[6] ,\c0|afi_addr[5] ,
\c0|afi_addr[4] ,\c0|afi_addr[3] ,\c0|afi_addr[2] ,\c0|afi_addr[1] ,\c0|afi_addr[0] }),
	.afi_ba({\c0|afi_ba[2] ,\c0|afi_ba[1] ,\c0|afi_ba[0] }),
	.afi_cke({\c0|afi_cke[1] ,\c0|afi_cke[0] }),
	.afi_cs_n({\c0|afi_cs_n[1] ,\c0|afi_cs_n[0] }),
	.afi_dm({\c0|afi_dm_int[9] ,\c0|afi_dm_int[8] ,\c0|afi_dm_int[7] ,\c0|afi_dm_int[6] ,\c0|afi_dm_int[5] ,\c0|afi_dm_int[4] ,\c0|afi_dm_int[3] ,\c0|afi_dm_int[2] ,\c0|afi_dm_int[1] ,\c0|afi_dm_int[0] }),
	.afi_dqs_burst({\c0|afi_dqs_burst[4] ,\c0|afi_dqs_burst[3] ,\c0|afi_dqs_burst[2] ,\c0|afi_dqs_burst[1] ,\c0|afi_dqs_burst[0] }),
	.afi_odt({\c0|afi_odt[1] ,\c0|afi_odt[0] }),
	.afi_rdata_en({\c0|afi_rdata_en[4] ,\c0|afi_rdata_en[3] ,\c0|afi_rdata_en[2] ,\c0|afi_rdata_en[1] ,\c0|afi_rdata_en[0] }),
	.afi_rdata_en_full({\c0|afi_rdata_en_full[4] ,\c0|afi_rdata_en_full[3] ,\c0|afi_rdata_en_full[2] ,\c0|afi_rdata_en_full[1] ,\c0|afi_rdata_en_full[0] }),
	.afi_wdata({\c0|afi_wdata_int[79] ,\c0|afi_wdata_int[78] ,\c0|afi_wdata_int[77] ,\c0|afi_wdata_int[76] ,\c0|afi_wdata_int[75] ,\c0|afi_wdata_int[74] ,\c0|afi_wdata_int[73] ,\c0|afi_wdata_int[72] ,\c0|afi_wdata_int[71] ,\c0|afi_wdata_int[70] ,\c0|afi_wdata_int[69] ,
\c0|afi_wdata_int[68] ,\c0|afi_wdata_int[67] ,\c0|afi_wdata_int[66] ,\c0|afi_wdata_int[65] ,\c0|afi_wdata_int[64] ,\c0|afi_wdata_int[63] ,\c0|afi_wdata_int[62] ,\c0|afi_wdata_int[61] ,\c0|afi_wdata_int[60] ,\c0|afi_wdata_int[59] ,\c0|afi_wdata_int[58] ,
\c0|afi_wdata_int[57] ,\c0|afi_wdata_int[56] ,\c0|afi_wdata_int[55] ,\c0|afi_wdata_int[54] ,\c0|afi_wdata_int[53] ,\c0|afi_wdata_int[52] ,\c0|afi_wdata_int[51] ,\c0|afi_wdata_int[50] ,\c0|afi_wdata_int[49] ,\c0|afi_wdata_int[48] ,\c0|afi_wdata_int[47] ,
\c0|afi_wdata_int[46] ,\c0|afi_wdata_int[45] ,\c0|afi_wdata_int[44] ,\c0|afi_wdata_int[43] ,\c0|afi_wdata_int[42] ,\c0|afi_wdata_int[41] ,\c0|afi_wdata_int[40] ,\c0|afi_wdata_int[39] ,\c0|afi_wdata_int[38] ,\c0|afi_wdata_int[37] ,\c0|afi_wdata_int[36] ,
\c0|afi_wdata_int[35] ,\c0|afi_wdata_int[34] ,\c0|afi_wdata_int[33] ,\c0|afi_wdata_int[32] ,\c0|afi_wdata_int[31] ,\c0|afi_wdata_int[30] ,\c0|afi_wdata_int[29] ,\c0|afi_wdata_int[28] ,\c0|afi_wdata_int[27] ,\c0|afi_wdata_int[26] ,\c0|afi_wdata_int[25] ,
\c0|afi_wdata_int[24] ,\c0|afi_wdata_int[23] ,\c0|afi_wdata_int[22] ,\c0|afi_wdata_int[21] ,\c0|afi_wdata_int[20] ,\c0|afi_wdata_int[19] ,\c0|afi_wdata_int[18] ,\c0|afi_wdata_int[17] ,\c0|afi_wdata_int[16] ,\c0|afi_wdata_int[15] ,\c0|afi_wdata_int[14] ,
\c0|afi_wdata_int[13] ,\c0|afi_wdata_int[12] ,\c0|afi_wdata_int[11] ,\c0|afi_wdata_int[10] ,\c0|afi_wdata_int[9] ,\c0|afi_wdata_int[8] ,\c0|afi_wdata_int[7] ,\c0|afi_wdata_int[6] ,\c0|afi_wdata_int[5] ,\c0|afi_wdata_int[4] ,\c0|afi_wdata_int[3] ,\c0|afi_wdata_int[2] ,
\c0|afi_wdata_int[1] ,\c0|afi_wdata_int[0] }),
	.afi_wdata_valid({\c0|afi_wdata_valid[4] ,\c0|afi_wdata_valid[3] ,\c0|afi_wdata_valid[2] ,\c0|afi_wdata_valid[1] ,\c0|afi_wdata_valid[0] }),
	.cfg_addlat({cfg_addlat_unconnected_wire_7,cfg_addlat_unconnected_wire_6,cfg_addlat_unconnected_wire_5,\c0|cfg_addlat_wire[4] ,\c0|cfg_addlat_wire[3] ,\c0|cfg_addlat_wire[2] ,\c0|cfg_addlat_wire[1] ,\c0|cfg_addlat_wire[0] }),
	.cfg_bankaddrwidth({cfg_bankaddrwidth_unconnected_wire_7,cfg_bankaddrwidth_unconnected_wire_6,cfg_bankaddrwidth_unconnected_wire_5,cfg_bankaddrwidth_unconnected_wire_4,cfg_bankaddrwidth_unconnected_wire_3,\c0|cfg_bankaddrwidth_wire[2] ,\c0|cfg_bankaddrwidth_wire[1] ,
\c0|cfg_bankaddrwidth_wire[0] }),
	.cfg_caswrlat({cfg_caswrlat_unconnected_wire_7,cfg_caswrlat_unconnected_wire_6,cfg_caswrlat_unconnected_wire_5,cfg_caswrlat_unconnected_wire_4,\c0|cfg_caswrlat_wire[3] ,\c0|cfg_caswrlat_wire[2] ,\c0|cfg_caswrlat_wire[1] ,\c0|cfg_caswrlat_wire[0] }),
	.cfg_coladdrwidth({cfg_coladdrwidth_unconnected_wire_7,cfg_coladdrwidth_unconnected_wire_6,cfg_coladdrwidth_unconnected_wire_5,\c0|cfg_coladdrwidth_wire[4] ,\c0|cfg_coladdrwidth_wire[3] ,\c0|cfg_coladdrwidth_wire[2] ,\c0|cfg_coladdrwidth_wire[1] ,\c0|cfg_coladdrwidth_wire[0] }),
	.cfg_csaddrwidth({cfg_csaddrwidth_unconnected_wire_7,cfg_csaddrwidth_unconnected_wire_6,cfg_csaddrwidth_unconnected_wire_5,cfg_csaddrwidth_unconnected_wire_4,cfg_csaddrwidth_unconnected_wire_3,\c0|cfg_csaddrwidth_wire[2] ,\c0|cfg_csaddrwidth_wire[1] ,\c0|cfg_csaddrwidth_wire[0] }),
	.cfg_devicewidth({cfg_devicewidth_unconnected_wire_7,cfg_devicewidth_unconnected_wire_6,cfg_devicewidth_unconnected_wire_5,cfg_devicewidth_unconnected_wire_4,\c0|cfg_devicewidth_wire[3] ,\c0|cfg_devicewidth_wire[2] ,\c0|cfg_devicewidth_wire[1] ,\c0|cfg_devicewidth_wire[0] }),
	.cfg_interfacewidth({\c0|cfg_interfacewidth_wire[7] ,\c0|cfg_interfacewidth_wire[6] ,\c0|cfg_interfacewidth_wire[5] ,\c0|cfg_interfacewidth_wire[4] ,\c0|cfg_interfacewidth_wire[3] ,\c0|cfg_interfacewidth_wire[2] ,\c0|cfg_interfacewidth_wire[1] ,\c0|cfg_interfacewidth_wire[0] }),
	.cfg_rowaddrwidth({cfg_rowaddrwidth_unconnected_wire_7,cfg_rowaddrwidth_unconnected_wire_6,cfg_rowaddrwidth_unconnected_wire_5,\c0|cfg_rowaddrwidth_wire[4] ,\c0|cfg_rowaddrwidth_wire[3] ,\c0|cfg_rowaddrwidth_wire[2] ,\c0|cfg_rowaddrwidth_wire[1] ,\c0|cfg_rowaddrwidth_wire[0] }),
	.cfg_tcl({cfg_tcl_unconnected_wire_7,cfg_tcl_unconnected_wire_6,cfg_tcl_unconnected_wire_5,\c0|cfg_tcl_wire[4] ,\c0|cfg_tcl_wire[3] ,\c0|cfg_tcl_wire[2] ,\c0|cfg_tcl_wire[1] ,\c0|cfg_tcl_wire[0] }),
	.cfg_tmrd({cfg_tmrd_unconnected_wire_7,cfg_tmrd_unconnected_wire_6,cfg_tmrd_unconnected_wire_5,cfg_tmrd_unconnected_wire_4,\c0|cfg_tmrd_wire[3] ,\c0|cfg_tmrd_wire[2] ,\c0|cfg_tmrd_wire[1] ,\c0|cfg_tmrd_wire[0] }),
	.cfg_trefi({cfg_trefi_unconnected_wire_15,cfg_trefi_unconnected_wire_14,cfg_trefi_unconnected_wire_13,\c0|cfg_trefi_wire[12] ,\c0|cfg_trefi_wire[11] ,\c0|cfg_trefi_wire[10] ,\c0|cfg_trefi_wire[9] ,\c0|cfg_trefi_wire[8] ,\c0|cfg_trefi_wire[7] ,\c0|cfg_trefi_wire[6] ,
\c0|cfg_trefi_wire[5] ,\c0|cfg_trefi_wire[4] ,\c0|cfg_trefi_wire[3] ,\c0|cfg_trefi_wire[2] ,\c0|cfg_trefi_wire[1] ,\c0|cfg_trefi_wire[0] }),
	.cfg_trfc({\c0|cfg_trfc_wire[7] ,\c0|cfg_trfc_wire[6] ,\c0|cfg_trfc_wire[5] ,\c0|cfg_trfc_wire[4] ,\c0|cfg_trfc_wire[3] ,\c0|cfg_trfc_wire[2] ,\c0|cfg_trfc_wire[1] ,\c0|cfg_trfc_wire[0] }),
	.cfg_twr({cfg_twr_unconnected_wire_7,cfg_twr_unconnected_wire_6,cfg_twr_unconnected_wire_5,cfg_twr_unconnected_wire_4,\c0|cfg_twr_wire[3] ,\c0|cfg_twr_wire[2] ,\c0|cfg_twr_wire[1] ,\c0|cfg_twr_wire[0] }),
	.afi_mem_clk_disable({\c0|afi_mem_clk_disable[0] }),
	.cfg_dramconfig({cfg_dramconfig_unconnected_wire_23,cfg_dramconfig_unconnected_wire_22,cfg_dramconfig_unconnected_wire_21,\c0|cfg_dramconfig_wire[20] ,\c0|cfg_dramconfig_wire[19] ,\c0|cfg_dramconfig_wire[18] ,\c0|cfg_dramconfig_wire[17] ,\c0|cfg_dramconfig_wire[16] ,
\c0|cfg_dramconfig_wire[15] ,\c0|cfg_dramconfig_wire[14] ,\c0|cfg_dramconfig_wire[13] ,\c0|cfg_dramconfig_wire[12] ,\c0|cfg_dramconfig_wire[11] ,\c0|cfg_dramconfig_wire[10] ,\c0|cfg_dramconfig_wire[9] ,\c0|cfg_dramconfig_wire[8] ,\c0|cfg_dramconfig_wire[7] ,
\c0|cfg_dramconfig_wire[6] ,\c0|cfg_dramconfig_wire[5] ,\c0|cfg_dramconfig_wire[4] ,\c0|cfg_dramconfig_wire[3] ,\c0|cfg_dramconfig_wire[2] ,\c0|cfg_dramconfig_wire[1] ,\c0|cfg_dramconfig_wire[0] }),
	.ctl_clk(\p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ));

Computer_System_hps_sdram_p0 p0(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(\pll|afi_clk ),
	.pll_write_clk(\pll|pll_write_clk ),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.afi_cal_fail(\p0|umemphy|afi_cal_fail ),
	.afi_cal_success(\p0|umemphy|afi_cal_success ),
	.afi_rdata_valid_0(\p0|umemphy|afi_rdata_valid[0] ),
	.ctl_reset_n(\p0|umemphy|ctl_reset_n ),
	.afi_rdata_0(\p0|umemphy|afi_rdata[0] ),
	.afi_rdata_1(\p0|umemphy|afi_rdata[1] ),
	.afi_rdata_2(\p0|umemphy|afi_rdata[2] ),
	.afi_rdata_3(\p0|umemphy|afi_rdata[3] ),
	.afi_rdata_4(\p0|umemphy|afi_rdata[4] ),
	.afi_rdata_5(\p0|umemphy|afi_rdata[5] ),
	.afi_rdata_6(\p0|umemphy|afi_rdata[6] ),
	.afi_rdata_7(\p0|umemphy|afi_rdata[7] ),
	.afi_rdata_8(\p0|umemphy|afi_rdata[8] ),
	.afi_rdata_9(\p0|umemphy|afi_rdata[9] ),
	.afi_rdata_10(\p0|umemphy|afi_rdata[10] ),
	.afi_rdata_11(\p0|umemphy|afi_rdata[11] ),
	.afi_rdata_12(\p0|umemphy|afi_rdata[12] ),
	.afi_rdata_13(\p0|umemphy|afi_rdata[13] ),
	.afi_rdata_14(\p0|umemphy|afi_rdata[14] ),
	.afi_rdata_15(\p0|umemphy|afi_rdata[15] ),
	.afi_rdata_16(\p0|umemphy|afi_rdata[16] ),
	.afi_rdata_17(\p0|umemphy|afi_rdata[17] ),
	.afi_rdata_18(\p0|umemphy|afi_rdata[18] ),
	.afi_rdata_19(\p0|umemphy|afi_rdata[19] ),
	.afi_rdata_20(\p0|umemphy|afi_rdata[20] ),
	.afi_rdata_21(\p0|umemphy|afi_rdata[21] ),
	.afi_rdata_22(\p0|umemphy|afi_rdata[22] ),
	.afi_rdata_23(\p0|umemphy|afi_rdata[23] ),
	.afi_rdata_24(\p0|umemphy|afi_rdata[24] ),
	.afi_rdata_25(\p0|umemphy|afi_rdata[25] ),
	.afi_rdata_26(\p0|umemphy|afi_rdata[26] ),
	.afi_rdata_27(\p0|umemphy|afi_rdata[27] ),
	.afi_rdata_28(\p0|umemphy|afi_rdata[28] ),
	.afi_rdata_29(\p0|umemphy|afi_rdata[29] ),
	.afi_rdata_30(\p0|umemphy|afi_rdata[30] ),
	.afi_rdata_31(\p0|umemphy|afi_rdata[31] ),
	.afi_rdata_32(\p0|umemphy|afi_rdata[32] ),
	.afi_rdata_33(\p0|umemphy|afi_rdata[33] ),
	.afi_rdata_34(\p0|umemphy|afi_rdata[34] ),
	.afi_rdata_35(\p0|umemphy|afi_rdata[35] ),
	.afi_rdata_36(\p0|umemphy|afi_rdata[36] ),
	.afi_rdata_37(\p0|umemphy|afi_rdata[37] ),
	.afi_rdata_38(\p0|umemphy|afi_rdata[38] ),
	.afi_rdata_39(\p0|umemphy|afi_rdata[39] ),
	.afi_rdata_40(\p0|umemphy|afi_rdata[40] ),
	.afi_rdata_41(\p0|umemphy|afi_rdata[41] ),
	.afi_rdata_42(\p0|umemphy|afi_rdata[42] ),
	.afi_rdata_43(\p0|umemphy|afi_rdata[43] ),
	.afi_rdata_44(\p0|umemphy|afi_rdata[44] ),
	.afi_rdata_45(\p0|umemphy|afi_rdata[45] ),
	.afi_rdata_46(\p0|umemphy|afi_rdata[46] ),
	.afi_rdata_47(\p0|umemphy|afi_rdata[47] ),
	.afi_rdata_48(\p0|umemphy|afi_rdata[48] ),
	.afi_rdata_49(\p0|umemphy|afi_rdata[49] ),
	.afi_rdata_50(\p0|umemphy|afi_rdata[50] ),
	.afi_rdata_51(\p0|umemphy|afi_rdata[51] ),
	.afi_rdata_52(\p0|umemphy|afi_rdata[52] ),
	.afi_rdata_53(\p0|umemphy|afi_rdata[53] ),
	.afi_rdata_54(\p0|umemphy|afi_rdata[54] ),
	.afi_rdata_55(\p0|umemphy|afi_rdata[55] ),
	.afi_rdata_56(\p0|umemphy|afi_rdata[56] ),
	.afi_rdata_57(\p0|umemphy|afi_rdata[57] ),
	.afi_rdata_58(\p0|umemphy|afi_rdata[58] ),
	.afi_rdata_59(\p0|umemphy|afi_rdata[59] ),
	.afi_rdata_60(\p0|umemphy|afi_rdata[60] ),
	.afi_rdata_61(\p0|umemphy|afi_rdata[61] ),
	.afi_rdata_62(\p0|umemphy|afi_rdata[62] ),
	.afi_rdata_63(\p0|umemphy|afi_rdata[63] ),
	.afi_rdata_64(\p0|umemphy|afi_rdata[64] ),
	.afi_rdata_65(\p0|umemphy|afi_rdata[65] ),
	.afi_rdata_66(\p0|umemphy|afi_rdata[66] ),
	.afi_rdata_67(\p0|umemphy|afi_rdata[67] ),
	.afi_rdata_68(\p0|umemphy|afi_rdata[68] ),
	.afi_rdata_69(\p0|umemphy|afi_rdata[69] ),
	.afi_rdata_70(\p0|umemphy|afi_rdata[70] ),
	.afi_rdata_71(\p0|umemphy|afi_rdata[71] ),
	.afi_rdata_72(\p0|umemphy|afi_rdata[72] ),
	.afi_rdata_73(\p0|umemphy|afi_rdata[73] ),
	.afi_rdata_74(\p0|umemphy|afi_rdata[74] ),
	.afi_rdata_75(\p0|umemphy|afi_rdata[75] ),
	.afi_rdata_76(\p0|umemphy|afi_rdata[76] ),
	.afi_rdata_77(\p0|umemphy|afi_rdata[77] ),
	.afi_rdata_78(\p0|umemphy|afi_rdata[78] ),
	.afi_rdata_79(\p0|umemphy|afi_rdata[79] ),
	.afi_wlat_0(\p0|umemphy|afi_wlat[0] ),
	.afi_wlat_1(\p0|umemphy|afi_wlat[1] ),
	.afi_wlat_2(\p0|umemphy|afi_wlat[2] ),
	.afi_wlat_3(\p0|umemphy|afi_wlat[3] ),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.afi_cas_n_0(\c0|afi_cas_n[0] ),
	.afi_ras_n_0(\c0|afi_ras_n[0] ),
	.afi_rst_n_0(\c0|afi_rst_n[0] ),
	.afi_we_n_0(\c0|afi_we_n[0] ),
	.afi_addr_0(\c0|afi_addr[0] ),
	.afi_addr_1(\c0|afi_addr[1] ),
	.afi_addr_2(\c0|afi_addr[2] ),
	.afi_addr_3(\c0|afi_addr[3] ),
	.afi_addr_4(\c0|afi_addr[4] ),
	.afi_addr_5(\c0|afi_addr[5] ),
	.afi_addr_6(\c0|afi_addr[6] ),
	.afi_addr_7(\c0|afi_addr[7] ),
	.afi_addr_8(\c0|afi_addr[8] ),
	.afi_addr_9(\c0|afi_addr[9] ),
	.afi_addr_10(\c0|afi_addr[10] ),
	.afi_addr_11(\c0|afi_addr[11] ),
	.afi_addr_12(\c0|afi_addr[12] ),
	.afi_addr_13(\c0|afi_addr[13] ),
	.afi_addr_14(\c0|afi_addr[14] ),
	.afi_addr_15(\c0|afi_addr[15] ),
	.afi_addr_16(\c0|afi_addr[16] ),
	.afi_addr_17(\c0|afi_addr[17] ),
	.afi_addr_18(\c0|afi_addr[18] ),
	.afi_addr_19(\c0|afi_addr[19] ),
	.afi_ba_0(\c0|afi_ba[0] ),
	.afi_ba_1(\c0|afi_ba[1] ),
	.afi_ba_2(\c0|afi_ba[2] ),
	.afi_cke_0(\c0|afi_cke[0] ),
	.afi_cke_1(\c0|afi_cke[1] ),
	.afi_cs_n_0(\c0|afi_cs_n[0] ),
	.afi_cs_n_1(\c0|afi_cs_n[1] ),
	.afi_dm_int_0(\c0|afi_dm_int[0] ),
	.afi_dm_int_1(\c0|afi_dm_int[1] ),
	.afi_dm_int_2(\c0|afi_dm_int[2] ),
	.afi_dm_int_3(\c0|afi_dm_int[3] ),
	.afi_dm_int_4(\c0|afi_dm_int[4] ),
	.afi_dm_int_5(\c0|afi_dm_int[5] ),
	.afi_dm_int_6(\c0|afi_dm_int[6] ),
	.afi_dm_int_7(\c0|afi_dm_int[7] ),
	.afi_dm_int_8(\c0|afi_dm_int[8] ),
	.afi_dm_int_9(\c0|afi_dm_int[9] ),
	.afi_dqs_burst_0(\c0|afi_dqs_burst[0] ),
	.afi_dqs_burst_1(\c0|afi_dqs_burst[1] ),
	.afi_dqs_burst_2(\c0|afi_dqs_burst[2] ),
	.afi_dqs_burst_3(\c0|afi_dqs_burst[3] ),
	.afi_dqs_burst_4(\c0|afi_dqs_burst[4] ),
	.afi_odt_0(\c0|afi_odt[0] ),
	.afi_odt_1(\c0|afi_odt[1] ),
	.afi_rdata_en_0(\c0|afi_rdata_en[0] ),
	.afi_rdata_en_1(\c0|afi_rdata_en[1] ),
	.afi_rdata_en_2(\c0|afi_rdata_en[2] ),
	.afi_rdata_en_3(\c0|afi_rdata_en[3] ),
	.afi_rdata_en_4(\c0|afi_rdata_en[4] ),
	.afi_rdata_en_full_0(\c0|afi_rdata_en_full[0] ),
	.afi_rdata_en_full_1(\c0|afi_rdata_en_full[1] ),
	.afi_rdata_en_full_2(\c0|afi_rdata_en_full[2] ),
	.afi_rdata_en_full_3(\c0|afi_rdata_en_full[3] ),
	.afi_rdata_en_full_4(\c0|afi_rdata_en_full[4] ),
	.afi_wdata_int_0(\c0|afi_wdata_int[0] ),
	.afi_wdata_int_1(\c0|afi_wdata_int[1] ),
	.afi_wdata_int_2(\c0|afi_wdata_int[2] ),
	.afi_wdata_int_3(\c0|afi_wdata_int[3] ),
	.afi_wdata_int_4(\c0|afi_wdata_int[4] ),
	.afi_wdata_int_5(\c0|afi_wdata_int[5] ),
	.afi_wdata_int_6(\c0|afi_wdata_int[6] ),
	.afi_wdata_int_7(\c0|afi_wdata_int[7] ),
	.afi_wdata_int_8(\c0|afi_wdata_int[8] ),
	.afi_wdata_int_9(\c0|afi_wdata_int[9] ),
	.afi_wdata_int_10(\c0|afi_wdata_int[10] ),
	.afi_wdata_int_11(\c0|afi_wdata_int[11] ),
	.afi_wdata_int_12(\c0|afi_wdata_int[12] ),
	.afi_wdata_int_13(\c0|afi_wdata_int[13] ),
	.afi_wdata_int_14(\c0|afi_wdata_int[14] ),
	.afi_wdata_int_15(\c0|afi_wdata_int[15] ),
	.afi_wdata_int_16(\c0|afi_wdata_int[16] ),
	.afi_wdata_int_17(\c0|afi_wdata_int[17] ),
	.afi_wdata_int_18(\c0|afi_wdata_int[18] ),
	.afi_wdata_int_19(\c0|afi_wdata_int[19] ),
	.afi_wdata_int_20(\c0|afi_wdata_int[20] ),
	.afi_wdata_int_21(\c0|afi_wdata_int[21] ),
	.afi_wdata_int_22(\c0|afi_wdata_int[22] ),
	.afi_wdata_int_23(\c0|afi_wdata_int[23] ),
	.afi_wdata_int_24(\c0|afi_wdata_int[24] ),
	.afi_wdata_int_25(\c0|afi_wdata_int[25] ),
	.afi_wdata_int_26(\c0|afi_wdata_int[26] ),
	.afi_wdata_int_27(\c0|afi_wdata_int[27] ),
	.afi_wdata_int_28(\c0|afi_wdata_int[28] ),
	.afi_wdata_int_29(\c0|afi_wdata_int[29] ),
	.afi_wdata_int_30(\c0|afi_wdata_int[30] ),
	.afi_wdata_int_31(\c0|afi_wdata_int[31] ),
	.afi_wdata_int_32(\c0|afi_wdata_int[32] ),
	.afi_wdata_int_33(\c0|afi_wdata_int[33] ),
	.afi_wdata_int_34(\c0|afi_wdata_int[34] ),
	.afi_wdata_int_35(\c0|afi_wdata_int[35] ),
	.afi_wdata_int_36(\c0|afi_wdata_int[36] ),
	.afi_wdata_int_37(\c0|afi_wdata_int[37] ),
	.afi_wdata_int_38(\c0|afi_wdata_int[38] ),
	.afi_wdata_int_39(\c0|afi_wdata_int[39] ),
	.afi_wdata_int_40(\c0|afi_wdata_int[40] ),
	.afi_wdata_int_41(\c0|afi_wdata_int[41] ),
	.afi_wdata_int_42(\c0|afi_wdata_int[42] ),
	.afi_wdata_int_43(\c0|afi_wdata_int[43] ),
	.afi_wdata_int_44(\c0|afi_wdata_int[44] ),
	.afi_wdata_int_45(\c0|afi_wdata_int[45] ),
	.afi_wdata_int_46(\c0|afi_wdata_int[46] ),
	.afi_wdata_int_47(\c0|afi_wdata_int[47] ),
	.afi_wdata_int_48(\c0|afi_wdata_int[48] ),
	.afi_wdata_int_49(\c0|afi_wdata_int[49] ),
	.afi_wdata_int_50(\c0|afi_wdata_int[50] ),
	.afi_wdata_int_51(\c0|afi_wdata_int[51] ),
	.afi_wdata_int_52(\c0|afi_wdata_int[52] ),
	.afi_wdata_int_53(\c0|afi_wdata_int[53] ),
	.afi_wdata_int_54(\c0|afi_wdata_int[54] ),
	.afi_wdata_int_55(\c0|afi_wdata_int[55] ),
	.afi_wdata_int_56(\c0|afi_wdata_int[56] ),
	.afi_wdata_int_57(\c0|afi_wdata_int[57] ),
	.afi_wdata_int_58(\c0|afi_wdata_int[58] ),
	.afi_wdata_int_59(\c0|afi_wdata_int[59] ),
	.afi_wdata_int_60(\c0|afi_wdata_int[60] ),
	.afi_wdata_int_61(\c0|afi_wdata_int[61] ),
	.afi_wdata_int_62(\c0|afi_wdata_int[62] ),
	.afi_wdata_int_63(\c0|afi_wdata_int[63] ),
	.afi_wdata_int_64(\c0|afi_wdata_int[64] ),
	.afi_wdata_int_65(\c0|afi_wdata_int[65] ),
	.afi_wdata_int_66(\c0|afi_wdata_int[66] ),
	.afi_wdata_int_67(\c0|afi_wdata_int[67] ),
	.afi_wdata_int_68(\c0|afi_wdata_int[68] ),
	.afi_wdata_int_69(\c0|afi_wdata_int[69] ),
	.afi_wdata_int_70(\c0|afi_wdata_int[70] ),
	.afi_wdata_int_71(\c0|afi_wdata_int[71] ),
	.afi_wdata_int_72(\c0|afi_wdata_int[72] ),
	.afi_wdata_int_73(\c0|afi_wdata_int[73] ),
	.afi_wdata_int_74(\c0|afi_wdata_int[74] ),
	.afi_wdata_int_75(\c0|afi_wdata_int[75] ),
	.afi_wdata_int_76(\c0|afi_wdata_int[76] ),
	.afi_wdata_int_77(\c0|afi_wdata_int[77] ),
	.afi_wdata_int_78(\c0|afi_wdata_int[78] ),
	.afi_wdata_int_79(\c0|afi_wdata_int[79] ),
	.afi_wdata_valid_0(\c0|afi_wdata_valid[0] ),
	.afi_wdata_valid_1(\c0|afi_wdata_valid[1] ),
	.afi_wdata_valid_2(\c0|afi_wdata_valid[2] ),
	.afi_wdata_valid_3(\c0|afi_wdata_valid[3] ),
	.afi_wdata_valid_4(\c0|afi_wdata_valid[4] ),
	.cfg_addlat_wire_0(\c0|cfg_addlat_wire[0] ),
	.cfg_addlat_wire_1(\c0|cfg_addlat_wire[1] ),
	.cfg_addlat_wire_2(\c0|cfg_addlat_wire[2] ),
	.cfg_addlat_wire_3(\c0|cfg_addlat_wire[3] ),
	.cfg_addlat_wire_4(\c0|cfg_addlat_wire[4] ),
	.cfg_bankaddrwidth_wire_0(\c0|cfg_bankaddrwidth_wire[0] ),
	.cfg_bankaddrwidth_wire_1(\c0|cfg_bankaddrwidth_wire[1] ),
	.cfg_bankaddrwidth_wire_2(\c0|cfg_bankaddrwidth_wire[2] ),
	.cfg_caswrlat_wire_0(\c0|cfg_caswrlat_wire[0] ),
	.cfg_caswrlat_wire_1(\c0|cfg_caswrlat_wire[1] ),
	.cfg_caswrlat_wire_2(\c0|cfg_caswrlat_wire[2] ),
	.cfg_caswrlat_wire_3(\c0|cfg_caswrlat_wire[3] ),
	.cfg_coladdrwidth_wire_0(\c0|cfg_coladdrwidth_wire[0] ),
	.cfg_coladdrwidth_wire_1(\c0|cfg_coladdrwidth_wire[1] ),
	.cfg_coladdrwidth_wire_2(\c0|cfg_coladdrwidth_wire[2] ),
	.cfg_coladdrwidth_wire_3(\c0|cfg_coladdrwidth_wire[3] ),
	.cfg_coladdrwidth_wire_4(\c0|cfg_coladdrwidth_wire[4] ),
	.cfg_csaddrwidth_wire_0(\c0|cfg_csaddrwidth_wire[0] ),
	.cfg_csaddrwidth_wire_1(\c0|cfg_csaddrwidth_wire[1] ),
	.cfg_csaddrwidth_wire_2(\c0|cfg_csaddrwidth_wire[2] ),
	.cfg_devicewidth_wire_0(\c0|cfg_devicewidth_wire[0] ),
	.cfg_devicewidth_wire_1(\c0|cfg_devicewidth_wire[1] ),
	.cfg_devicewidth_wire_2(\c0|cfg_devicewidth_wire[2] ),
	.cfg_devicewidth_wire_3(\c0|cfg_devicewidth_wire[3] ),
	.cfg_interfacewidth_wire_0(\c0|cfg_interfacewidth_wire[0] ),
	.cfg_interfacewidth_wire_1(\c0|cfg_interfacewidth_wire[1] ),
	.cfg_interfacewidth_wire_2(\c0|cfg_interfacewidth_wire[2] ),
	.cfg_interfacewidth_wire_3(\c0|cfg_interfacewidth_wire[3] ),
	.cfg_interfacewidth_wire_4(\c0|cfg_interfacewidth_wire[4] ),
	.cfg_interfacewidth_wire_5(\c0|cfg_interfacewidth_wire[5] ),
	.cfg_interfacewidth_wire_6(\c0|cfg_interfacewidth_wire[6] ),
	.cfg_interfacewidth_wire_7(\c0|cfg_interfacewidth_wire[7] ),
	.cfg_rowaddrwidth_wire_0(\c0|cfg_rowaddrwidth_wire[0] ),
	.cfg_rowaddrwidth_wire_1(\c0|cfg_rowaddrwidth_wire[1] ),
	.cfg_rowaddrwidth_wire_2(\c0|cfg_rowaddrwidth_wire[2] ),
	.cfg_rowaddrwidth_wire_3(\c0|cfg_rowaddrwidth_wire[3] ),
	.cfg_rowaddrwidth_wire_4(\c0|cfg_rowaddrwidth_wire[4] ),
	.cfg_tcl_wire_0(\c0|cfg_tcl_wire[0] ),
	.cfg_tcl_wire_1(\c0|cfg_tcl_wire[1] ),
	.cfg_tcl_wire_2(\c0|cfg_tcl_wire[2] ),
	.cfg_tcl_wire_3(\c0|cfg_tcl_wire[3] ),
	.cfg_tcl_wire_4(\c0|cfg_tcl_wire[4] ),
	.cfg_tmrd_wire_0(\c0|cfg_tmrd_wire[0] ),
	.cfg_tmrd_wire_1(\c0|cfg_tmrd_wire[1] ),
	.cfg_tmrd_wire_2(\c0|cfg_tmrd_wire[2] ),
	.cfg_tmrd_wire_3(\c0|cfg_tmrd_wire[3] ),
	.cfg_trefi_wire_0(\c0|cfg_trefi_wire[0] ),
	.cfg_trefi_wire_1(\c0|cfg_trefi_wire[1] ),
	.cfg_trefi_wire_2(\c0|cfg_trefi_wire[2] ),
	.cfg_trefi_wire_3(\c0|cfg_trefi_wire[3] ),
	.cfg_trefi_wire_4(\c0|cfg_trefi_wire[4] ),
	.cfg_trefi_wire_5(\c0|cfg_trefi_wire[5] ),
	.cfg_trefi_wire_6(\c0|cfg_trefi_wire[6] ),
	.cfg_trefi_wire_7(\c0|cfg_trefi_wire[7] ),
	.cfg_trefi_wire_8(\c0|cfg_trefi_wire[8] ),
	.cfg_trefi_wire_9(\c0|cfg_trefi_wire[9] ),
	.cfg_trefi_wire_10(\c0|cfg_trefi_wire[10] ),
	.cfg_trefi_wire_11(\c0|cfg_trefi_wire[11] ),
	.cfg_trefi_wire_12(\c0|cfg_trefi_wire[12] ),
	.cfg_trfc_wire_0(\c0|cfg_trfc_wire[0] ),
	.cfg_trfc_wire_1(\c0|cfg_trfc_wire[1] ),
	.cfg_trfc_wire_2(\c0|cfg_trfc_wire[2] ),
	.cfg_trfc_wire_3(\c0|cfg_trfc_wire[3] ),
	.cfg_trfc_wire_4(\c0|cfg_trfc_wire[4] ),
	.cfg_trfc_wire_5(\c0|cfg_trfc_wire[5] ),
	.cfg_trfc_wire_6(\c0|cfg_trfc_wire[6] ),
	.cfg_trfc_wire_7(\c0|cfg_trfc_wire[7] ),
	.cfg_twr_wire_0(\c0|cfg_twr_wire[0] ),
	.cfg_twr_wire_1(\c0|cfg_twr_wire[1] ),
	.cfg_twr_wire_2(\c0|cfg_twr_wire[2] ),
	.cfg_twr_wire_3(\c0|cfg_twr_wire[3] ),
	.afi_mem_clk_disable_0(\c0|afi_mem_clk_disable[0] ),
	.cfg_dramconfig_wire_0(\c0|cfg_dramconfig_wire[0] ),
	.cfg_dramconfig_wire_1(\c0|cfg_dramconfig_wire[1] ),
	.cfg_dramconfig_wire_2(\c0|cfg_dramconfig_wire[2] ),
	.cfg_dramconfig_wire_3(\c0|cfg_dramconfig_wire[3] ),
	.cfg_dramconfig_wire_4(\c0|cfg_dramconfig_wire[4] ),
	.cfg_dramconfig_wire_5(\c0|cfg_dramconfig_wire[5] ),
	.cfg_dramconfig_wire_6(\c0|cfg_dramconfig_wire[6] ),
	.cfg_dramconfig_wire_7(\c0|cfg_dramconfig_wire[7] ),
	.cfg_dramconfig_wire_8(\c0|cfg_dramconfig_wire[8] ),
	.cfg_dramconfig_wire_9(\c0|cfg_dramconfig_wire[9] ),
	.cfg_dramconfig_wire_10(\c0|cfg_dramconfig_wire[10] ),
	.cfg_dramconfig_wire_11(\c0|cfg_dramconfig_wire[11] ),
	.cfg_dramconfig_wire_12(\c0|cfg_dramconfig_wire[12] ),
	.cfg_dramconfig_wire_13(\c0|cfg_dramconfig_wire[13] ),
	.cfg_dramconfig_wire_14(\c0|cfg_dramconfig_wire[14] ),
	.cfg_dramconfig_wire_15(\c0|cfg_dramconfig_wire[15] ),
	.cfg_dramconfig_wire_16(\c0|cfg_dramconfig_wire[16] ),
	.cfg_dramconfig_wire_17(\c0|cfg_dramconfig_wire[17] ),
	.cfg_dramconfig_wire_18(\c0|cfg_dramconfig_wire[18] ),
	.cfg_dramconfig_wire_19(\c0|cfg_dramconfig_wire[19] ),
	.cfg_dramconfig_wire_20(\c0|cfg_dramconfig_wire[20] ),
	.ctl_clk(\p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ),
	.dll_delayctrl_0(\dll|dll_delayctrl[0] ),
	.dll_delayctrl_1(\dll|dll_delayctrl[1] ),
	.dll_delayctrl_2(\dll|dll_delayctrl[2] ),
	.dll_delayctrl_3(\dll|dll_delayctrl[3] ),
	.dll_delayctrl_4(\dll|dll_delayctrl[4] ),
	.dll_delayctrl_5(\dll|dll_delayctrl[5] ),
	.dll_delayctrl_6(\dll|dll_delayctrl[6] ),
	.GND_port(GND_port));

Computer_System_hps_sdram_pll pll(
	.pll_mem_clk(\pll|afi_clk ),
	.pll_write_clk(\pll|pll_write_clk ));

endmodule

module Computer_System_altera_mem_if_dll_cyclonev (
	clk,
	dll_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	clk;
output 	[6:0] dll_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [6:0] dll_wys_m_DELAYCTRLOUT_bus;

assign dll_delayctrl[0] = dll_wys_m_DELAYCTRLOUT_bus[0];
assign dll_delayctrl[1] = dll_wys_m_DELAYCTRLOUT_bus[1];
assign dll_delayctrl[2] = dll_wys_m_DELAYCTRLOUT_bus[2];
assign dll_delayctrl[3] = dll_wys_m_DELAYCTRLOUT_bus[3];
assign dll_delayctrl[4] = dll_wys_m_DELAYCTRLOUT_bus[4];
assign dll_delayctrl[5] = dll_wys_m_DELAYCTRLOUT_bus[5];
assign dll_delayctrl[6] = dll_wys_m_DELAYCTRLOUT_bus[6];

cyclonev_dll dll_wys_m(
	.clk(clk),
	.aload(vcc),
	.upndnin(gnd),
	.upndninclkena(gnd),
	.dqsupdate(),
	.upndnout(),
	.delayctrlout(dll_wys_m_DELAYCTRLOUT_bus));
defparam dll_wys_m.delayctrlout_mode = "normal";
defparam dll_wys_m.input_frequency = "2500 ps";
defparam dll_wys_m.jitter_reduction = "true";
defparam dll_wys_m.sim_buffer_delay_increment = 10;
defparam dll_wys_m.sim_buffer_intrinsic_delay = 175;
defparam dll_wys_m.sim_valid_lock = 16;
defparam dll_wys_m.sim_valid_lockcount = 0;
defparam dll_wys_m.static_delay_ctrl = 8;
defparam dll_wys_m.upndnout_mode = "clock";
defparam dll_wys_m.use_upndnin = "false";
defparam dll_wys_m.use_upndninclkena = "false";

endmodule

module Computer_System_altera_mem_if_hard_memory_controller_top_cyclonev (
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid,
	ctl_reset_n,
	afi_rdata,
	afi_wlat,
	afi_cas_n,
	afi_ras_n,
	afi_rst_n,
	afi_we_n,
	afi_addr,
	afi_ba,
	afi_cke,
	afi_cs_n,
	afi_dm,
	afi_dqs_burst,
	afi_odt,
	afi_rdata_en,
	afi_rdata_en_full,
	afi_wdata,
	afi_wdata_valid,
	cfg_addlat,
	cfg_bankaddrwidth,
	cfg_caswrlat,
	cfg_coladdrwidth,
	cfg_csaddrwidth,
	cfg_devicewidth,
	cfg_interfacewidth,
	cfg_rowaddrwidth,
	cfg_tcl,
	cfg_tmrd,
	cfg_trefi,
	cfg_trfc,
	cfg_twr,
	afi_mem_clk_disable,
	cfg_dramconfig,
	ctl_clk)/* synthesis synthesis_greybox=0 */;
input 	afi_cal_fail;
input 	afi_cal_success;
input 	[0:0] afi_rdata_valid;
input 	ctl_reset_n;
input 	[79:0] afi_rdata;
input 	[3:0] afi_wlat;
output 	[0:0] afi_cas_n;
output 	[0:0] afi_ras_n;
output 	[0:0] afi_rst_n;
output 	[0:0] afi_we_n;
output 	[19:0] afi_addr;
output 	[2:0] afi_ba;
output 	[1:0] afi_cke;
output 	[1:0] afi_cs_n;
output 	[9:0] afi_dm;
output 	[4:0] afi_dqs_burst;
output 	[1:0] afi_odt;
output 	[4:0] afi_rdata_en;
output 	[4:0] afi_rdata_en_full;
output 	[79:0] afi_wdata;
output 	[4:0] afi_wdata_valid;
output 	[7:0] cfg_addlat;
output 	[7:0] cfg_bankaddrwidth;
output 	[7:0] cfg_caswrlat;
output 	[7:0] cfg_coladdrwidth;
output 	[7:0] cfg_csaddrwidth;
output 	[7:0] cfg_devicewidth;
output 	[7:0] cfg_interfacewidth;
output 	[7:0] cfg_rowaddrwidth;
output 	[7:0] cfg_tcl;
output 	[7:0] cfg_tmrd;
output 	[15:0] cfg_trefi;
output 	[7:0] cfg_trfc;
output 	[7:0] cfg_twr;
output 	[0:0] afi_mem_clk_disable;
output 	[23:0] cfg_dramconfig;
input 	ctl_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [19:0] hmc_inst_AFIADDR_bus;
wire [2:0] hmc_inst_AFIBA_bus;
wire [1:0] hmc_inst_AFICKE_bus;
wire [1:0] hmc_inst_AFICSN_bus;
wire [9:0] hmc_inst_AFIDM_bus;
wire [4:0] hmc_inst_AFIDQSBURST_bus;
wire [1:0] hmc_inst_AFIODT_bus;
wire [4:0] hmc_inst_AFIRDATAEN_bus;
wire [4:0] hmc_inst_AFIRDATAENFULL_bus;
wire [79:0] hmc_inst_AFIWDATA_bus;
wire [4:0] hmc_inst_AFIWDATAVALID_bus;
wire [4:0] hmc_inst_CFGADDLAT_bus;
wire [2:0] hmc_inst_CFGBANKADDRWIDTH_bus;
wire [3:0] hmc_inst_CFGCASWRLAT_bus;
wire [4:0] hmc_inst_CFGCOLADDRWIDTH_bus;
wire [2:0] hmc_inst_CFGCSADDRWIDTH_bus;
wire [3:0] hmc_inst_CFGDEVICEWIDTH_bus;
wire [7:0] hmc_inst_CFGINTERFACEWIDTH_bus;
wire [4:0] hmc_inst_CFGROWADDRWIDTH_bus;
wire [4:0] hmc_inst_CFGTCL_bus;
wire [3:0] hmc_inst_CFGTMRD_bus;
wire [12:0] hmc_inst_CFGTREFI_bus;
wire [7:0] hmc_inst_CFGTRFC_bus;
wire [3:0] hmc_inst_CFGTWR_bus;
wire [1:0] hmc_inst_CTLMEMCLKDISABLE_bus;
wire [20:0] hmc_inst_DRAMCONFIG_bus;

assign afi_addr[0] = hmc_inst_AFIADDR_bus[0];
assign afi_addr[1] = hmc_inst_AFIADDR_bus[1];
assign afi_addr[2] = hmc_inst_AFIADDR_bus[2];
assign afi_addr[3] = hmc_inst_AFIADDR_bus[3];
assign afi_addr[4] = hmc_inst_AFIADDR_bus[4];
assign afi_addr[5] = hmc_inst_AFIADDR_bus[5];
assign afi_addr[6] = hmc_inst_AFIADDR_bus[6];
assign afi_addr[7] = hmc_inst_AFIADDR_bus[7];
assign afi_addr[8] = hmc_inst_AFIADDR_bus[8];
assign afi_addr[9] = hmc_inst_AFIADDR_bus[9];
assign afi_addr[10] = hmc_inst_AFIADDR_bus[10];
assign afi_addr[11] = hmc_inst_AFIADDR_bus[11];
assign afi_addr[12] = hmc_inst_AFIADDR_bus[12];
assign afi_addr[13] = hmc_inst_AFIADDR_bus[13];
assign afi_addr[14] = hmc_inst_AFIADDR_bus[14];
assign afi_addr[15] = hmc_inst_AFIADDR_bus[15];
assign afi_addr[16] = hmc_inst_AFIADDR_bus[16];
assign afi_addr[17] = hmc_inst_AFIADDR_bus[17];
assign afi_addr[18] = hmc_inst_AFIADDR_bus[18];
assign afi_addr[19] = hmc_inst_AFIADDR_bus[19];

assign afi_ba[0] = hmc_inst_AFIBA_bus[0];
assign afi_ba[1] = hmc_inst_AFIBA_bus[1];
assign afi_ba[2] = hmc_inst_AFIBA_bus[2];

assign afi_cke[0] = hmc_inst_AFICKE_bus[0];
assign afi_cke[1] = hmc_inst_AFICKE_bus[1];

assign afi_cs_n[0] = hmc_inst_AFICSN_bus[0];
assign afi_cs_n[1] = hmc_inst_AFICSN_bus[1];

assign afi_dm[0] = hmc_inst_AFIDM_bus[0];
assign afi_dm[1] = hmc_inst_AFIDM_bus[1];
assign afi_dm[2] = hmc_inst_AFIDM_bus[2];
assign afi_dm[3] = hmc_inst_AFIDM_bus[3];
assign afi_dm[4] = hmc_inst_AFIDM_bus[4];
assign afi_dm[5] = hmc_inst_AFIDM_bus[5];
assign afi_dm[6] = hmc_inst_AFIDM_bus[6];
assign afi_dm[7] = hmc_inst_AFIDM_bus[7];
assign afi_dm[8] = hmc_inst_AFIDM_bus[8];
assign afi_dm[9] = hmc_inst_AFIDM_bus[9];

assign afi_dqs_burst[0] = hmc_inst_AFIDQSBURST_bus[0];
assign afi_dqs_burst[1] = hmc_inst_AFIDQSBURST_bus[1];
assign afi_dqs_burst[2] = hmc_inst_AFIDQSBURST_bus[2];
assign afi_dqs_burst[3] = hmc_inst_AFIDQSBURST_bus[3];
assign afi_dqs_burst[4] = hmc_inst_AFIDQSBURST_bus[4];

assign afi_odt[0] = hmc_inst_AFIODT_bus[0];
assign afi_odt[1] = hmc_inst_AFIODT_bus[1];

assign afi_rdata_en[0] = hmc_inst_AFIRDATAEN_bus[0];
assign afi_rdata_en[1] = hmc_inst_AFIRDATAEN_bus[1];
assign afi_rdata_en[2] = hmc_inst_AFIRDATAEN_bus[2];
assign afi_rdata_en[3] = hmc_inst_AFIRDATAEN_bus[3];
assign afi_rdata_en[4] = hmc_inst_AFIRDATAEN_bus[4];

assign afi_rdata_en_full[0] = hmc_inst_AFIRDATAENFULL_bus[0];
assign afi_rdata_en_full[1] = hmc_inst_AFIRDATAENFULL_bus[1];
assign afi_rdata_en_full[2] = hmc_inst_AFIRDATAENFULL_bus[2];
assign afi_rdata_en_full[3] = hmc_inst_AFIRDATAENFULL_bus[3];
assign afi_rdata_en_full[4] = hmc_inst_AFIRDATAENFULL_bus[4];

assign afi_wdata[0] = hmc_inst_AFIWDATA_bus[0];
assign afi_wdata[1] = hmc_inst_AFIWDATA_bus[1];
assign afi_wdata[2] = hmc_inst_AFIWDATA_bus[2];
assign afi_wdata[3] = hmc_inst_AFIWDATA_bus[3];
assign afi_wdata[4] = hmc_inst_AFIWDATA_bus[4];
assign afi_wdata[5] = hmc_inst_AFIWDATA_bus[5];
assign afi_wdata[6] = hmc_inst_AFIWDATA_bus[6];
assign afi_wdata[7] = hmc_inst_AFIWDATA_bus[7];
assign afi_wdata[8] = hmc_inst_AFIWDATA_bus[8];
assign afi_wdata[9] = hmc_inst_AFIWDATA_bus[9];
assign afi_wdata[10] = hmc_inst_AFIWDATA_bus[10];
assign afi_wdata[11] = hmc_inst_AFIWDATA_bus[11];
assign afi_wdata[12] = hmc_inst_AFIWDATA_bus[12];
assign afi_wdata[13] = hmc_inst_AFIWDATA_bus[13];
assign afi_wdata[14] = hmc_inst_AFIWDATA_bus[14];
assign afi_wdata[15] = hmc_inst_AFIWDATA_bus[15];
assign afi_wdata[16] = hmc_inst_AFIWDATA_bus[16];
assign afi_wdata[17] = hmc_inst_AFIWDATA_bus[17];
assign afi_wdata[18] = hmc_inst_AFIWDATA_bus[18];
assign afi_wdata[19] = hmc_inst_AFIWDATA_bus[19];
assign afi_wdata[20] = hmc_inst_AFIWDATA_bus[20];
assign afi_wdata[21] = hmc_inst_AFIWDATA_bus[21];
assign afi_wdata[22] = hmc_inst_AFIWDATA_bus[22];
assign afi_wdata[23] = hmc_inst_AFIWDATA_bus[23];
assign afi_wdata[24] = hmc_inst_AFIWDATA_bus[24];
assign afi_wdata[25] = hmc_inst_AFIWDATA_bus[25];
assign afi_wdata[26] = hmc_inst_AFIWDATA_bus[26];
assign afi_wdata[27] = hmc_inst_AFIWDATA_bus[27];
assign afi_wdata[28] = hmc_inst_AFIWDATA_bus[28];
assign afi_wdata[29] = hmc_inst_AFIWDATA_bus[29];
assign afi_wdata[30] = hmc_inst_AFIWDATA_bus[30];
assign afi_wdata[31] = hmc_inst_AFIWDATA_bus[31];
assign afi_wdata[32] = hmc_inst_AFIWDATA_bus[32];
assign afi_wdata[33] = hmc_inst_AFIWDATA_bus[33];
assign afi_wdata[34] = hmc_inst_AFIWDATA_bus[34];
assign afi_wdata[35] = hmc_inst_AFIWDATA_bus[35];
assign afi_wdata[36] = hmc_inst_AFIWDATA_bus[36];
assign afi_wdata[37] = hmc_inst_AFIWDATA_bus[37];
assign afi_wdata[38] = hmc_inst_AFIWDATA_bus[38];
assign afi_wdata[39] = hmc_inst_AFIWDATA_bus[39];
assign afi_wdata[40] = hmc_inst_AFIWDATA_bus[40];
assign afi_wdata[41] = hmc_inst_AFIWDATA_bus[41];
assign afi_wdata[42] = hmc_inst_AFIWDATA_bus[42];
assign afi_wdata[43] = hmc_inst_AFIWDATA_bus[43];
assign afi_wdata[44] = hmc_inst_AFIWDATA_bus[44];
assign afi_wdata[45] = hmc_inst_AFIWDATA_bus[45];
assign afi_wdata[46] = hmc_inst_AFIWDATA_bus[46];
assign afi_wdata[47] = hmc_inst_AFIWDATA_bus[47];
assign afi_wdata[48] = hmc_inst_AFIWDATA_bus[48];
assign afi_wdata[49] = hmc_inst_AFIWDATA_bus[49];
assign afi_wdata[50] = hmc_inst_AFIWDATA_bus[50];
assign afi_wdata[51] = hmc_inst_AFIWDATA_bus[51];
assign afi_wdata[52] = hmc_inst_AFIWDATA_bus[52];
assign afi_wdata[53] = hmc_inst_AFIWDATA_bus[53];
assign afi_wdata[54] = hmc_inst_AFIWDATA_bus[54];
assign afi_wdata[55] = hmc_inst_AFIWDATA_bus[55];
assign afi_wdata[56] = hmc_inst_AFIWDATA_bus[56];
assign afi_wdata[57] = hmc_inst_AFIWDATA_bus[57];
assign afi_wdata[58] = hmc_inst_AFIWDATA_bus[58];
assign afi_wdata[59] = hmc_inst_AFIWDATA_bus[59];
assign afi_wdata[60] = hmc_inst_AFIWDATA_bus[60];
assign afi_wdata[61] = hmc_inst_AFIWDATA_bus[61];
assign afi_wdata[62] = hmc_inst_AFIWDATA_bus[62];
assign afi_wdata[63] = hmc_inst_AFIWDATA_bus[63];
assign afi_wdata[64] = hmc_inst_AFIWDATA_bus[64];
assign afi_wdata[65] = hmc_inst_AFIWDATA_bus[65];
assign afi_wdata[66] = hmc_inst_AFIWDATA_bus[66];
assign afi_wdata[67] = hmc_inst_AFIWDATA_bus[67];
assign afi_wdata[68] = hmc_inst_AFIWDATA_bus[68];
assign afi_wdata[69] = hmc_inst_AFIWDATA_bus[69];
assign afi_wdata[70] = hmc_inst_AFIWDATA_bus[70];
assign afi_wdata[71] = hmc_inst_AFIWDATA_bus[71];
assign afi_wdata[72] = hmc_inst_AFIWDATA_bus[72];
assign afi_wdata[73] = hmc_inst_AFIWDATA_bus[73];
assign afi_wdata[74] = hmc_inst_AFIWDATA_bus[74];
assign afi_wdata[75] = hmc_inst_AFIWDATA_bus[75];
assign afi_wdata[76] = hmc_inst_AFIWDATA_bus[76];
assign afi_wdata[77] = hmc_inst_AFIWDATA_bus[77];
assign afi_wdata[78] = hmc_inst_AFIWDATA_bus[78];
assign afi_wdata[79] = hmc_inst_AFIWDATA_bus[79];

assign afi_wdata_valid[0] = hmc_inst_AFIWDATAVALID_bus[0];
assign afi_wdata_valid[1] = hmc_inst_AFIWDATAVALID_bus[1];
assign afi_wdata_valid[2] = hmc_inst_AFIWDATAVALID_bus[2];
assign afi_wdata_valid[3] = hmc_inst_AFIWDATAVALID_bus[3];
assign afi_wdata_valid[4] = hmc_inst_AFIWDATAVALID_bus[4];

assign cfg_addlat[0] = hmc_inst_CFGADDLAT_bus[0];
assign cfg_addlat[1] = hmc_inst_CFGADDLAT_bus[1];
assign cfg_addlat[2] = hmc_inst_CFGADDLAT_bus[2];
assign cfg_addlat[3] = hmc_inst_CFGADDLAT_bus[3];
assign cfg_addlat[4] = hmc_inst_CFGADDLAT_bus[4];

assign cfg_bankaddrwidth[0] = hmc_inst_CFGBANKADDRWIDTH_bus[0];
assign cfg_bankaddrwidth[1] = hmc_inst_CFGBANKADDRWIDTH_bus[1];
assign cfg_bankaddrwidth[2] = hmc_inst_CFGBANKADDRWIDTH_bus[2];

assign cfg_caswrlat[0] = hmc_inst_CFGCASWRLAT_bus[0];
assign cfg_caswrlat[1] = hmc_inst_CFGCASWRLAT_bus[1];
assign cfg_caswrlat[2] = hmc_inst_CFGCASWRLAT_bus[2];
assign cfg_caswrlat[3] = hmc_inst_CFGCASWRLAT_bus[3];

assign cfg_coladdrwidth[0] = hmc_inst_CFGCOLADDRWIDTH_bus[0];
assign cfg_coladdrwidth[1] = hmc_inst_CFGCOLADDRWIDTH_bus[1];
assign cfg_coladdrwidth[2] = hmc_inst_CFGCOLADDRWIDTH_bus[2];
assign cfg_coladdrwidth[3] = hmc_inst_CFGCOLADDRWIDTH_bus[3];
assign cfg_coladdrwidth[4] = hmc_inst_CFGCOLADDRWIDTH_bus[4];

assign cfg_csaddrwidth[0] = hmc_inst_CFGCSADDRWIDTH_bus[0];
assign cfg_csaddrwidth[1] = hmc_inst_CFGCSADDRWIDTH_bus[1];
assign cfg_csaddrwidth[2] = hmc_inst_CFGCSADDRWIDTH_bus[2];

assign cfg_devicewidth[0] = hmc_inst_CFGDEVICEWIDTH_bus[0];
assign cfg_devicewidth[1] = hmc_inst_CFGDEVICEWIDTH_bus[1];
assign cfg_devicewidth[2] = hmc_inst_CFGDEVICEWIDTH_bus[2];
assign cfg_devicewidth[3] = hmc_inst_CFGDEVICEWIDTH_bus[3];

assign cfg_interfacewidth[0] = hmc_inst_CFGINTERFACEWIDTH_bus[0];
assign cfg_interfacewidth[1] = hmc_inst_CFGINTERFACEWIDTH_bus[1];
assign cfg_interfacewidth[2] = hmc_inst_CFGINTERFACEWIDTH_bus[2];
assign cfg_interfacewidth[3] = hmc_inst_CFGINTERFACEWIDTH_bus[3];
assign cfg_interfacewidth[4] = hmc_inst_CFGINTERFACEWIDTH_bus[4];
assign cfg_interfacewidth[5] = hmc_inst_CFGINTERFACEWIDTH_bus[5];
assign cfg_interfacewidth[6] = hmc_inst_CFGINTERFACEWIDTH_bus[6];
assign cfg_interfacewidth[7] = hmc_inst_CFGINTERFACEWIDTH_bus[7];

assign cfg_rowaddrwidth[0] = hmc_inst_CFGROWADDRWIDTH_bus[0];
assign cfg_rowaddrwidth[1] = hmc_inst_CFGROWADDRWIDTH_bus[1];
assign cfg_rowaddrwidth[2] = hmc_inst_CFGROWADDRWIDTH_bus[2];
assign cfg_rowaddrwidth[3] = hmc_inst_CFGROWADDRWIDTH_bus[3];
assign cfg_rowaddrwidth[4] = hmc_inst_CFGROWADDRWIDTH_bus[4];

assign cfg_tcl[0] = hmc_inst_CFGTCL_bus[0];
assign cfg_tcl[1] = hmc_inst_CFGTCL_bus[1];
assign cfg_tcl[2] = hmc_inst_CFGTCL_bus[2];
assign cfg_tcl[3] = hmc_inst_CFGTCL_bus[3];
assign cfg_tcl[4] = hmc_inst_CFGTCL_bus[4];

assign cfg_tmrd[0] = hmc_inst_CFGTMRD_bus[0];
assign cfg_tmrd[1] = hmc_inst_CFGTMRD_bus[1];
assign cfg_tmrd[2] = hmc_inst_CFGTMRD_bus[2];
assign cfg_tmrd[3] = hmc_inst_CFGTMRD_bus[3];

assign cfg_trefi[0] = hmc_inst_CFGTREFI_bus[0];
assign cfg_trefi[1] = hmc_inst_CFGTREFI_bus[1];
assign cfg_trefi[2] = hmc_inst_CFGTREFI_bus[2];
assign cfg_trefi[3] = hmc_inst_CFGTREFI_bus[3];
assign cfg_trefi[4] = hmc_inst_CFGTREFI_bus[4];
assign cfg_trefi[5] = hmc_inst_CFGTREFI_bus[5];
assign cfg_trefi[6] = hmc_inst_CFGTREFI_bus[6];
assign cfg_trefi[7] = hmc_inst_CFGTREFI_bus[7];
assign cfg_trefi[8] = hmc_inst_CFGTREFI_bus[8];
assign cfg_trefi[9] = hmc_inst_CFGTREFI_bus[9];
assign cfg_trefi[10] = hmc_inst_CFGTREFI_bus[10];
assign cfg_trefi[11] = hmc_inst_CFGTREFI_bus[11];
assign cfg_trefi[12] = hmc_inst_CFGTREFI_bus[12];

assign cfg_trfc[0] = hmc_inst_CFGTRFC_bus[0];
assign cfg_trfc[1] = hmc_inst_CFGTRFC_bus[1];
assign cfg_trfc[2] = hmc_inst_CFGTRFC_bus[2];
assign cfg_trfc[3] = hmc_inst_CFGTRFC_bus[3];
assign cfg_trfc[4] = hmc_inst_CFGTRFC_bus[4];
assign cfg_trfc[5] = hmc_inst_CFGTRFC_bus[5];
assign cfg_trfc[6] = hmc_inst_CFGTRFC_bus[6];
assign cfg_trfc[7] = hmc_inst_CFGTRFC_bus[7];

assign cfg_twr[0] = hmc_inst_CFGTWR_bus[0];
assign cfg_twr[1] = hmc_inst_CFGTWR_bus[1];
assign cfg_twr[2] = hmc_inst_CFGTWR_bus[2];
assign cfg_twr[3] = hmc_inst_CFGTWR_bus[3];

assign afi_mem_clk_disable[0] = hmc_inst_CTLMEMCLKDISABLE_bus[0];

assign cfg_dramconfig[0] = hmc_inst_DRAMCONFIG_bus[0];
assign cfg_dramconfig[1] = hmc_inst_DRAMCONFIG_bus[1];
assign cfg_dramconfig[2] = hmc_inst_DRAMCONFIG_bus[2];
assign cfg_dramconfig[3] = hmc_inst_DRAMCONFIG_bus[3];
assign cfg_dramconfig[4] = hmc_inst_DRAMCONFIG_bus[4];
assign cfg_dramconfig[5] = hmc_inst_DRAMCONFIG_bus[5];
assign cfg_dramconfig[6] = hmc_inst_DRAMCONFIG_bus[6];
assign cfg_dramconfig[7] = hmc_inst_DRAMCONFIG_bus[7];
assign cfg_dramconfig[8] = hmc_inst_DRAMCONFIG_bus[8];
assign cfg_dramconfig[9] = hmc_inst_DRAMCONFIG_bus[9];
assign cfg_dramconfig[10] = hmc_inst_DRAMCONFIG_bus[10];
assign cfg_dramconfig[11] = hmc_inst_DRAMCONFIG_bus[11];
assign cfg_dramconfig[12] = hmc_inst_DRAMCONFIG_bus[12];
assign cfg_dramconfig[13] = hmc_inst_DRAMCONFIG_bus[13];
assign cfg_dramconfig[14] = hmc_inst_DRAMCONFIG_bus[14];
assign cfg_dramconfig[15] = hmc_inst_DRAMCONFIG_bus[15];
assign cfg_dramconfig[16] = hmc_inst_DRAMCONFIG_bus[16];
assign cfg_dramconfig[17] = hmc_inst_DRAMCONFIG_bus[17];
assign cfg_dramconfig[18] = hmc_inst_DRAMCONFIG_bus[18];
assign cfg_dramconfig[19] = hmc_inst_DRAMCONFIG_bus[19];
assign cfg_dramconfig[20] = hmc_inst_DRAMCONFIG_bus[20];

cyclonev_hmc hmc_inst(
	.afirdatavalid(afi_rdata_valid[0]),
	.csrclk(gnd),
	.csrdin(gnd),
	.csren(gnd),
	.ctlcalfail(afi_cal_fail),
	.ctlcalsuccess(afi_cal_success),
	.ctlclk(ctl_clk),
	.ctlresetn(ctl_reset_n),
	.globalresetn(gnd),
	.iavstcmdresetn0(vcc),
	.iavstcmdresetn1(vcc),
	.iavstcmdresetn2(vcc),
	.iavstcmdresetn3(vcc),
	.iavstcmdresetn4(vcc),
	.iavstcmdresetn5(vcc),
	.iavstrdclk0(gnd),
	.iavstrdclk1(gnd),
	.iavstrdclk2(gnd),
	.iavstrdclk3(gnd),
	.iavstrdready0(vcc),
	.iavstrdready1(vcc),
	.iavstrdready2(vcc),
	.iavstrdready3(vcc),
	.iavstrdresetn0(vcc),
	.iavstrdresetn1(vcc),
	.iavstrdresetn2(vcc),
	.iavstrdresetn3(vcc),
	.iavstwrackready0(vcc),
	.iavstwrackready1(vcc),
	.iavstwrackready2(vcc),
	.iavstwrackready3(vcc),
	.iavstwrackready4(vcc),
	.iavstwrackready5(vcc),
	.iavstwrclk0(gnd),
	.iavstwrclk1(gnd),
	.iavstwrclk2(gnd),
	.iavstwrclk3(gnd),
	.iavstwrresetn0(vcc),
	.iavstwrresetn1(vcc),
	.iavstwrresetn2(vcc),
	.iavstwrresetn3(vcc),
	.localdeeppowerdnreq(gnd),
	.localrefreshreq(gnd),
	.localselfrfshreq(gnd),
	.mmrbe(gnd),
	.mmrburstbegin(vcc),
	.mmrclk(gnd),
	.mmrreadreq(gnd),
	.mmrresetn(vcc),
	.mmrwritereq(gnd),
	.portclk0(gnd),
	.portclk1(gnd),
	.portclk2(gnd),
	.portclk3(gnd),
	.portclk4(gnd),
	.portclk5(gnd),
	.scanenable(gnd),
	.scbe(gnd),
	.scburstbegin(gnd),
	.scclk(gnd),
	.screadreq(gnd),
	.scresetn(vcc),
	.scwritereq(gnd),
	.afirdata({afi_rdata[79],afi_rdata[78],afi_rdata[77],afi_rdata[76],afi_rdata[75],afi_rdata[74],afi_rdata[73],afi_rdata[72],afi_rdata[71],afi_rdata[70],afi_rdata[69],afi_rdata[68],afi_rdata[67],afi_rdata[66],afi_rdata[65],afi_rdata[64],afi_rdata[63],afi_rdata[62],afi_rdata[61],afi_rdata[60],afi_rdata[59],afi_rdata[58],afi_rdata[57],afi_rdata[56],afi_rdata[55],afi_rdata[54],afi_rdata[53],afi_rdata[52],
afi_rdata[51],afi_rdata[50],afi_rdata[49],afi_rdata[48],afi_rdata[47],afi_rdata[46],afi_rdata[45],afi_rdata[44],afi_rdata[43],afi_rdata[42],afi_rdata[41],afi_rdata[40],afi_rdata[39],afi_rdata[38],afi_rdata[37],afi_rdata[36],afi_rdata[35],afi_rdata[34],afi_rdata[33],afi_rdata[32],afi_rdata[31],afi_rdata[30],afi_rdata[29],afi_rdata[28],afi_rdata[27],afi_rdata[26],afi_rdata[25],afi_rdata[24],
afi_rdata[23],afi_rdata[22],afi_rdata[21],afi_rdata[20],afi_rdata[19],afi_rdata[18],afi_rdata[17],afi_rdata[16],afi_rdata[15],afi_rdata[14],afi_rdata[13],afi_rdata[12],afi_rdata[11],afi_rdata[10],afi_rdata[9],afi_rdata[8],afi_rdata[7],afi_rdata[6],afi_rdata[5],afi_rdata[4],afi_rdata[3],afi_rdata[2],afi_rdata[1],afi_rdata[0]}),
	.afiseqbusy({gnd,gnd}),
	.afiwlat({afi_wlat[3],afi_wlat[2],afi_wlat[1],afi_wlat[0]}),
	.bondingin1({gnd,gnd,gnd,gnd}),
	.bondingin2({gnd,gnd,gnd,gnd,gnd,gnd}),
	.bondingin3({gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata0({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata1({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata2({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata3({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata4({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata5({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata0({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata1({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata2({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata3({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.localdeeppowerdnchip({gnd,gnd}),
	.localrefreshchip({gnd,gnd}),
	.localselfrfshchip({gnd,gnd}),
	.mmraddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.mmrburstcount({gnd,vcc}),
	.mmrwdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.scaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.scburstcount({gnd,gnd}),
	.scwdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.aficasn(afi_cas_n[0]),
	.afirasn(afi_ras_n[0]),
	.afirstn(afi_rst_n[0]),
	.afiwen(afi_we_n[0]),
	.csrdout(),
	.ctlcalreq(),
	.ctlinitreq(),
	.localdeeppowerdnack(),
	.localinitdone(),
	.localpowerdownack(),
	.localrefreshack(),
	.localselfrfshack(),
	.localstsctlempty(),
	.mmrrdatavalid(),
	.mmrwaitrequest(),
	.oammready0(),
	.oammready1(),
	.oammready2(),
	.oammready3(),
	.oammready4(),
	.oammready5(),
	.ordavstvalid0(),
	.ordavstvalid1(),
	.ordavstvalid2(),
	.ordavstvalid3(),
	.owrackavstdata0(),
	.owrackavstdata1(),
	.owrackavstdata2(),
	.owrackavstdata3(),
	.owrackavstdata4(),
	.owrackavstdata5(),
	.owrackavstvalid0(),
	.owrackavstvalid1(),
	.owrackavstvalid2(),
	.owrackavstvalid3(),
	.owrackavstvalid4(),
	.owrackavstvalid5(),
	.scrdatavalid(),
	.scwaitrequest(),
	.afiaddr(hmc_inst_AFIADDR_bus),
	.afiba(hmc_inst_AFIBA_bus),
	.aficke(hmc_inst_AFICKE_bus),
	.aficsn(hmc_inst_AFICSN_bus),
	.afictllongidle(),
	.afictlrefreshdone(),
	.afidm(hmc_inst_AFIDM_bus),
	.afidqsburst(hmc_inst_AFIDQSBURST_bus),
	.afiodt(hmc_inst_AFIODT_bus),
	.afirdataen(hmc_inst_AFIRDATAEN_bus),
	.afirdataenfull(hmc_inst_AFIRDATAENFULL_bus),
	.afiwdata(hmc_inst_AFIWDATA_bus),
	.afiwdatavalid(hmc_inst_AFIWDATAVALID_bus),
	.bondingout1(),
	.bondingout2(),
	.bondingout3(),
	.cfgaddlat(hmc_inst_CFGADDLAT_bus),
	.cfgbankaddrwidth(hmc_inst_CFGBANKADDRWIDTH_bus),
	.cfgcaswrlat(hmc_inst_CFGCASWRLAT_bus),
	.cfgcoladdrwidth(hmc_inst_CFGCOLADDRWIDTH_bus),
	.cfgcsaddrwidth(hmc_inst_CFGCSADDRWIDTH_bus),
	.cfgdevicewidth(hmc_inst_CFGDEVICEWIDTH_bus),
	.cfginterfacewidth(hmc_inst_CFGINTERFACEWIDTH_bus),
	.cfgrowaddrwidth(hmc_inst_CFGROWADDRWIDTH_bus),
	.cfgtcl(hmc_inst_CFGTCL_bus),
	.cfgtmrd(hmc_inst_CFGTMRD_bus),
	.cfgtrefi(hmc_inst_CFGTREFI_bus),
	.cfgtrfc(hmc_inst_CFGTRFC_bus),
	.cfgtwr(hmc_inst_CFGTWR_bus),
	.ctlcalbytelaneseln(),
	.ctlmemclkdisable(hmc_inst_CTLMEMCLKDISABLE_bus),
	.dramconfig(hmc_inst_DRAMCONFIG_bus),
	.mmrrdata(),
	.ordavstdata0(),
	.ordavstdata1(),
	.ordavstdata2(),
	.ordavstdata3(),
	.scrdata());
defparam hmc_inst.attr_counter_one_mask = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_one_match = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_one_reset = "disabled";
defparam hmc_inst.attr_counter_zero_mask = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_zero_match = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_zero_reset = "disabled";
defparam hmc_inst.attr_debug_select_byte = 32'b00000000000000000000000000000000;
defparam hmc_inst.attr_static_config_valid = "disabled";
defparam hmc_inst.auto_pch_enable_0 = "disabled";
defparam hmc_inst.auto_pch_enable_1 = "disabled";
defparam hmc_inst.auto_pch_enable_2 = "disabled";
defparam hmc_inst.auto_pch_enable_3 = "disabled";
defparam hmc_inst.auto_pch_enable_4 = "disabled";
defparam hmc_inst.auto_pch_enable_5 = "disabled";
defparam hmc_inst.cal_req = "disabled";
defparam hmc_inst.cfg_burst_length = "bl_8";
defparam hmc_inst.cfg_interface_width = "dwidth_32";
defparam hmc_inst.cfg_self_rfsh_exit_cycles = "self_rfsh_exit_cycles_512";
defparam hmc_inst.cfg_starve_limit = "starve_limit_10";
defparam hmc_inst.cfg_type = "ddr3";
defparam hmc_inst.clr_intr = "no_clr_intr";
defparam hmc_inst.cmd_port_in_use_0 = "false";
defparam hmc_inst.cmd_port_in_use_1 = "false";
defparam hmc_inst.cmd_port_in_use_2 = "false";
defparam hmc_inst.cmd_port_in_use_3 = "false";
defparam hmc_inst.cmd_port_in_use_4 = "false";
defparam hmc_inst.cmd_port_in_use_5 = "false";
defparam hmc_inst.cport0_rdy_almost_full = "not_full";
defparam hmc_inst.cport0_rfifo_map = "fifo_0";
defparam hmc_inst.cport0_type = "disable";
defparam hmc_inst.cport0_wfifo_map = "fifo_0";
defparam hmc_inst.cport1_rdy_almost_full = "not_full";
defparam hmc_inst.cport1_rfifo_map = "fifo_0";
defparam hmc_inst.cport1_type = "disable";
defparam hmc_inst.cport1_wfifo_map = "fifo_0";
defparam hmc_inst.cport2_rdy_almost_full = "not_full";
defparam hmc_inst.cport2_rfifo_map = "fifo_0";
defparam hmc_inst.cport2_type = "disable";
defparam hmc_inst.cport2_wfifo_map = "fifo_0";
defparam hmc_inst.cport3_rdy_almost_full = "not_full";
defparam hmc_inst.cport3_rfifo_map = "fifo_0";
defparam hmc_inst.cport3_type = "disable";
defparam hmc_inst.cport3_wfifo_map = "fifo_0";
defparam hmc_inst.cport4_rdy_almost_full = "not_full";
defparam hmc_inst.cport4_rfifo_map = "fifo_0";
defparam hmc_inst.cport4_type = "disable";
defparam hmc_inst.cport4_wfifo_map = "fifo_0";
defparam hmc_inst.cport5_rdy_almost_full = "not_full";
defparam hmc_inst.cport5_rfifo_map = "fifo_0";
defparam hmc_inst.cport5_type = "disable";
defparam hmc_inst.cport5_wfifo_map = "fifo_0";
defparam hmc_inst.ctl_addr_order = "chip_row_bank_col";
defparam hmc_inst.ctl_ecc_enabled = "ctl_ecc_disabled";
defparam hmc_inst.ctl_ecc_rmw_enabled = "ctl_ecc_rmw_disabled";
defparam hmc_inst.ctl_regdimm_enabled = "regdimm_disabled";
defparam hmc_inst.ctl_usr_refresh = "ctl_usr_refresh_disabled";
defparam hmc_inst.ctrl_width = "data_width_64_bit";
defparam hmc_inst.cyc_to_rld_jars_0 = 1;
defparam hmc_inst.cyc_to_rld_jars_1 = 1;
defparam hmc_inst.cyc_to_rld_jars_2 = 1;
defparam hmc_inst.cyc_to_rld_jars_3 = 1;
defparam hmc_inst.cyc_to_rld_jars_4 = 1;
defparam hmc_inst.cyc_to_rld_jars_5 = 1;
defparam hmc_inst.delay_bonding = "bonding_latency_0";
defparam hmc_inst.dfx_bypass_enable = "dfx_bypass_disabled";
defparam hmc_inst.disable_merging = "merging_enabled";
defparam hmc_inst.ecc_dq_width = "ecc_dq_width_0";
defparam hmc_inst.enable_atpg = "disabled";
defparam hmc_inst.enable_bonding_0 = "disabled";
defparam hmc_inst.enable_bonding_1 = "disabled";
defparam hmc_inst.enable_bonding_2 = "disabled";
defparam hmc_inst.enable_bonding_3 = "disabled";
defparam hmc_inst.enable_bonding_4 = "disabled";
defparam hmc_inst.enable_bonding_5 = "disabled";
defparam hmc_inst.enable_bonding_wrapback = "disabled";
defparam hmc_inst.enable_burst_interrupt = "disabled";
defparam hmc_inst.enable_burst_terminate = "disabled";
defparam hmc_inst.enable_dqs_tracking = "enabled";
defparam hmc_inst.enable_ecc_code_overwrites = "disabled";
defparam hmc_inst.enable_fast_exit_ppd = "disabled";
defparam hmc_inst.enable_intr = "disabled";
defparam hmc_inst.enable_no_dm = "disabled";
defparam hmc_inst.enable_pipelineglobal = "disabled";
defparam hmc_inst.extra_ctl_clk_act_to_act = 0;
defparam hmc_inst.extra_ctl_clk_act_to_act_diff_bank = 0;
defparam hmc_inst.extra_ctl_clk_act_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_act_to_rdwr = 0;
defparam hmc_inst.extra_ctl_clk_arf_period = 0;
defparam hmc_inst.extra_ctl_clk_arf_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_four_act_to_act = 0;
defparam hmc_inst.extra_ctl_clk_pch_all_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_pch_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_pdn_period = 0;
defparam hmc_inst.extra_ctl_clk_pdn_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_rd_ap_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_rd = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_rd_diff_chip = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_wr = 2;
defparam hmc_inst.extra_ctl_clk_rd_to_wr_bc = 2;
defparam hmc_inst.extra_ctl_clk_rd_to_wr_diff_chip = 2;
defparam hmc_inst.extra_ctl_clk_srf_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_srf_to_zq_cal = 0;
defparam hmc_inst.extra_ctl_clk_wr_ap_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_rd = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_rd_bc = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_rd_diff_chip = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_wr = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_wr_diff_chip = 0;
defparam hmc_inst.gen_dbe = "gen_dbe_disabled";
defparam hmc_inst.gen_sbe = "gen_sbe_disabled";
defparam hmc_inst.inc_sync = "fifo_set_2";
defparam hmc_inst.local_if_cs_width = "addr_width_0";
defparam hmc_inst.mask_corr_dropped_intr = "disabled";
defparam hmc_inst.mask_dbe_intr = "disabled";
defparam hmc_inst.mask_sbe_intr = "disabled";
defparam hmc_inst.mem_auto_pd_cycles = 0;
defparam hmc_inst.mem_clk_entry_cycles = 10;
defparam hmc_inst.mem_if_al = "al_0";
defparam hmc_inst.mem_if_bankaddr_width = "addr_width_3";
defparam hmc_inst.mem_if_burstlength = "mem_if_burstlength_8";
defparam hmc_inst.mem_if_coladdr_width = "addr_width_10";
defparam hmc_inst.mem_if_cs_per_rank = "mem_if_cs_per_rank_1";
defparam hmc_inst.mem_if_cs_width = "mem_if_cs_width_1";
defparam hmc_inst.mem_if_dq_per_chip = "mem_if_dq_per_chip_8";
defparam hmc_inst.mem_if_dqs_width = "dqs_width_4";
defparam hmc_inst.mem_if_dwidth = "mem_if_dwidth_32";
defparam hmc_inst.mem_if_memtype = "ddr3_sdram";
defparam hmc_inst.mem_if_rowaddr_width = "addr_width_15";
defparam hmc_inst.mem_if_speedbin = "ddr3_1600_8_8_8";
defparam hmc_inst.mem_if_tccd = "tccd_4";
defparam hmc_inst.mem_if_tcl = "tcl_11";
defparam hmc_inst.mem_if_tcwl = "tcwl_8";
defparam hmc_inst.mem_if_tfaw = "tfaw_12";
defparam hmc_inst.mem_if_tmrd = "tmrd_4";
defparam hmc_inst.mem_if_tras = "tras_14";
defparam hmc_inst.mem_if_trc = "trc_20";
defparam hmc_inst.mem_if_trcd = "trcd_6";
defparam hmc_inst.mem_if_trefi = 3120;
defparam hmc_inst.mem_if_trfc = 104;
defparam hmc_inst.mem_if_trp = "trp_6";
defparam hmc_inst.mem_if_trrd = "trrd_3";
defparam hmc_inst.mem_if_trtp = "trtp_3";
defparam hmc_inst.mem_if_twr = "twr_6";
defparam hmc_inst.mem_if_twtr = "twtr_4";
defparam hmc_inst.mmr_cfg_mem_bl = "mp_bl_8";
defparam hmc_inst.output_regd = "disabled";
defparam hmc_inst.pdn_exit_cycles = "slow_exit";
defparam hmc_inst.port0_width = "port_32_bit";
defparam hmc_inst.port1_width = "port_32_bit";
defparam hmc_inst.port2_width = "port_32_bit";
defparam hmc_inst.port3_width = "port_32_bit";
defparam hmc_inst.port4_width = "port_32_bit";
defparam hmc_inst.port5_width = "port_32_bit";
defparam hmc_inst.power_saving_exit_cycles = 5;
defparam hmc_inst.priority_0_0 = "weight_0";
defparam hmc_inst.priority_0_1 = "weight_0";
defparam hmc_inst.priority_0_2 = "weight_0";
defparam hmc_inst.priority_0_3 = "weight_0";
defparam hmc_inst.priority_0_4 = "weight_0";
defparam hmc_inst.priority_0_5 = "weight_0";
defparam hmc_inst.priority_1_0 = "weight_0";
defparam hmc_inst.priority_1_1 = "weight_0";
defparam hmc_inst.priority_1_2 = "weight_0";
defparam hmc_inst.priority_1_3 = "weight_0";
defparam hmc_inst.priority_1_4 = "weight_0";
defparam hmc_inst.priority_1_5 = "weight_0";
defparam hmc_inst.priority_2_0 = "weight_0";
defparam hmc_inst.priority_2_1 = "weight_0";
defparam hmc_inst.priority_2_2 = "weight_0";
defparam hmc_inst.priority_2_3 = "weight_0";
defparam hmc_inst.priority_2_4 = "weight_0";
defparam hmc_inst.priority_2_5 = "weight_0";
defparam hmc_inst.priority_3_0 = "weight_0";
defparam hmc_inst.priority_3_1 = "weight_0";
defparam hmc_inst.priority_3_2 = "weight_0";
defparam hmc_inst.priority_3_3 = "weight_0";
defparam hmc_inst.priority_3_4 = "weight_0";
defparam hmc_inst.priority_3_5 = "weight_0";
defparam hmc_inst.priority_4_0 = "weight_0";
defparam hmc_inst.priority_4_1 = "weight_0";
defparam hmc_inst.priority_4_2 = "weight_0";
defparam hmc_inst.priority_4_3 = "weight_0";
defparam hmc_inst.priority_4_4 = "weight_0";
defparam hmc_inst.priority_4_5 = "weight_0";
defparam hmc_inst.priority_5_0 = "weight_0";
defparam hmc_inst.priority_5_1 = "weight_0";
defparam hmc_inst.priority_5_2 = "weight_0";
defparam hmc_inst.priority_5_3 = "weight_0";
defparam hmc_inst.priority_5_4 = "weight_0";
defparam hmc_inst.priority_5_5 = "weight_0";
defparam hmc_inst.priority_6_0 = "weight_0";
defparam hmc_inst.priority_6_1 = "weight_0";
defparam hmc_inst.priority_6_2 = "weight_0";
defparam hmc_inst.priority_6_3 = "weight_0";
defparam hmc_inst.priority_6_4 = "weight_0";
defparam hmc_inst.priority_6_5 = "weight_0";
defparam hmc_inst.priority_7_0 = "weight_0";
defparam hmc_inst.priority_7_1 = "weight_0";
defparam hmc_inst.priority_7_2 = "weight_0";
defparam hmc_inst.priority_7_3 = "weight_0";
defparam hmc_inst.priority_7_4 = "weight_0";
defparam hmc_inst.priority_7_5 = "weight_0";
defparam hmc_inst.priority_remap = 0;
defparam hmc_inst.rcfg_static_weight_0 = "weight_0";
defparam hmc_inst.rcfg_static_weight_1 = "weight_0";
defparam hmc_inst.rcfg_static_weight_2 = "weight_0";
defparam hmc_inst.rcfg_static_weight_3 = "weight_0";
defparam hmc_inst.rcfg_static_weight_4 = "weight_0";
defparam hmc_inst.rcfg_static_weight_5 = "weight_0";
defparam hmc_inst.rcfg_sum_wt_priority_0 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_1 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_2 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_3 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_4 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_5 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_6 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_7 = 0;
defparam hmc_inst.rcfg_user_priority_0 = "priority_1";
defparam hmc_inst.rcfg_user_priority_1 = "priority_1";
defparam hmc_inst.rcfg_user_priority_2 = "priority_1";
defparam hmc_inst.rcfg_user_priority_3 = "priority_1";
defparam hmc_inst.rcfg_user_priority_4 = "priority_1";
defparam hmc_inst.rcfg_user_priority_5 = "priority_1";
defparam hmc_inst.rd_dwidth_0 = "dwidth_0";
defparam hmc_inst.rd_dwidth_1 = "dwidth_0";
defparam hmc_inst.rd_dwidth_2 = "dwidth_0";
defparam hmc_inst.rd_dwidth_3 = "dwidth_0";
defparam hmc_inst.rd_dwidth_4 = "dwidth_0";
defparam hmc_inst.rd_dwidth_5 = "dwidth_0";
defparam hmc_inst.rd_fifo_in_use_0 = "false";
defparam hmc_inst.rd_fifo_in_use_1 = "false";
defparam hmc_inst.rd_fifo_in_use_2 = "false";
defparam hmc_inst.rd_fifo_in_use_3 = "false";
defparam hmc_inst.rd_port_info_0 = "use_no";
defparam hmc_inst.rd_port_info_1 = "use_no";
defparam hmc_inst.rd_port_info_2 = "use_no";
defparam hmc_inst.rd_port_info_3 = "use_no";
defparam hmc_inst.rd_port_info_4 = "use_no";
defparam hmc_inst.rd_port_info_5 = "use_no";
defparam hmc_inst.read_odt_chip = "odt_disabled";
defparam hmc_inst.reorder_data = "data_reordering";
defparam hmc_inst.rfifo0_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo1_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo2_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo3_cport_map = "cmd_port_0";
defparam hmc_inst.single_ready_0 = "concatenate_rdy";
defparam hmc_inst.single_ready_1 = "concatenate_rdy";
defparam hmc_inst.single_ready_2 = "concatenate_rdy";
defparam hmc_inst.single_ready_3 = "concatenate_rdy";
defparam hmc_inst.static_weight_0 = "weight_0";
defparam hmc_inst.static_weight_1 = "weight_0";
defparam hmc_inst.static_weight_2 = "weight_0";
defparam hmc_inst.static_weight_3 = "weight_0";
defparam hmc_inst.static_weight_4 = "weight_0";
defparam hmc_inst.static_weight_5 = "weight_0";
defparam hmc_inst.sum_wt_priority_0 = 0;
defparam hmc_inst.sum_wt_priority_1 = 0;
defparam hmc_inst.sum_wt_priority_2 = 0;
defparam hmc_inst.sum_wt_priority_3 = 0;
defparam hmc_inst.sum_wt_priority_4 = 0;
defparam hmc_inst.sum_wt_priority_5 = 0;
defparam hmc_inst.sum_wt_priority_6 = 0;
defparam hmc_inst.sum_wt_priority_7 = 0;
defparam hmc_inst.sync_mode_0 = "asynchronous";
defparam hmc_inst.sync_mode_1 = "asynchronous";
defparam hmc_inst.sync_mode_2 = "asynchronous";
defparam hmc_inst.sync_mode_3 = "asynchronous";
defparam hmc_inst.sync_mode_4 = "asynchronous";
defparam hmc_inst.sync_mode_5 = "asynchronous";
defparam hmc_inst.test_mode = "normal_mode";
defparam hmc_inst.thld_jar1_0 = "threshold_32";
defparam hmc_inst.thld_jar1_1 = "threshold_32";
defparam hmc_inst.thld_jar1_2 = "threshold_32";
defparam hmc_inst.thld_jar1_3 = "threshold_32";
defparam hmc_inst.thld_jar1_4 = "threshold_32";
defparam hmc_inst.thld_jar1_5 = "threshold_32";
defparam hmc_inst.thld_jar2_0 = "threshold_16";
defparam hmc_inst.thld_jar2_1 = "threshold_16";
defparam hmc_inst.thld_jar2_2 = "threshold_16";
defparam hmc_inst.thld_jar2_3 = "threshold_16";
defparam hmc_inst.thld_jar2_4 = "threshold_16";
defparam hmc_inst.thld_jar2_5 = "threshold_16";
defparam hmc_inst.use_almost_empty_0 = "empty";
defparam hmc_inst.use_almost_empty_1 = "empty";
defparam hmc_inst.use_almost_empty_2 = "empty";
defparam hmc_inst.use_almost_empty_3 = "empty";
defparam hmc_inst.user_ecc_en = "disable";
defparam hmc_inst.user_priority_0 = "priority_1";
defparam hmc_inst.user_priority_1 = "priority_1";
defparam hmc_inst.user_priority_2 = "priority_1";
defparam hmc_inst.user_priority_3 = "priority_1";
defparam hmc_inst.user_priority_4 = "priority_1";
defparam hmc_inst.user_priority_5 = "priority_1";
defparam hmc_inst.wfifo0_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo0_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo1_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo1_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo2_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo2_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo3_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo3_rdy_almost_full = "not_full";
defparam hmc_inst.wr_dwidth_0 = "dwidth_0";
defparam hmc_inst.wr_dwidth_1 = "dwidth_0";
defparam hmc_inst.wr_dwidth_2 = "dwidth_0";
defparam hmc_inst.wr_dwidth_3 = "dwidth_0";
defparam hmc_inst.wr_dwidth_4 = "dwidth_0";
defparam hmc_inst.wr_dwidth_5 = "dwidth_0";
defparam hmc_inst.wr_fifo_in_use_0 = "false";
defparam hmc_inst.wr_fifo_in_use_1 = "false";
defparam hmc_inst.wr_fifo_in_use_2 = "false";
defparam hmc_inst.wr_fifo_in_use_3 = "false";
defparam hmc_inst.wr_port_info_0 = "use_no";
defparam hmc_inst.wr_port_info_1 = "use_no";
defparam hmc_inst.wr_port_info_2 = "use_no";
defparam hmc_inst.wr_port_info_3 = "use_no";
defparam hmc_inst.wr_port_info_4 = "use_no";
defparam hmc_inst.wr_port_info_5 = "use_no";
defparam hmc_inst.write_odt_chip = "write_chip0_odt0_chip1";

endmodule

module Computer_System_altera_mem_if_oct_cyclonev (
	parallelterminationcontrol,
	seriesterminationcontrol,
	oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	[15:0] parallelterminationcontrol;
output 	[15:0] seriesterminationcontrol;
input 	oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sd1a_0~O_CLKUSRDFTOUT ;
wire \wire_sd1a_serdataout[0] ;

wire [15:0] sd2a_0_PARALLELTERMINATIONCONTROL_bus;
wire [15:0] sd2a_0_SERIESTERMINATIONCONTROL_bus;

assign parallelterminationcontrol[0] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[0];
assign parallelterminationcontrol[1] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[1];
assign parallelterminationcontrol[2] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[2];
assign parallelterminationcontrol[3] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[3];
assign parallelterminationcontrol[4] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[4];
assign parallelterminationcontrol[5] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[5];
assign parallelterminationcontrol[6] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[6];
assign parallelterminationcontrol[7] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[7];
assign parallelterminationcontrol[8] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[8];
assign parallelterminationcontrol[9] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[9];
assign parallelterminationcontrol[10] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[10];
assign parallelterminationcontrol[11] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[11];
assign parallelterminationcontrol[12] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[12];
assign parallelterminationcontrol[13] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[13];
assign parallelterminationcontrol[14] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[14];
assign parallelterminationcontrol[15] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[15];

assign seriesterminationcontrol[0] = sd2a_0_SERIESTERMINATIONCONTROL_bus[0];
assign seriesterminationcontrol[1] = sd2a_0_SERIESTERMINATIONCONTROL_bus[1];
assign seriesterminationcontrol[2] = sd2a_0_SERIESTERMINATIONCONTROL_bus[2];
assign seriesterminationcontrol[3] = sd2a_0_SERIESTERMINATIONCONTROL_bus[3];
assign seriesterminationcontrol[4] = sd2a_0_SERIESTERMINATIONCONTROL_bus[4];
assign seriesterminationcontrol[5] = sd2a_0_SERIESTERMINATIONCONTROL_bus[5];
assign seriesterminationcontrol[6] = sd2a_0_SERIESTERMINATIONCONTROL_bus[6];
assign seriesterminationcontrol[7] = sd2a_0_SERIESTERMINATIONCONTROL_bus[7];
assign seriesterminationcontrol[8] = sd2a_0_SERIESTERMINATIONCONTROL_bus[8];
assign seriesterminationcontrol[9] = sd2a_0_SERIESTERMINATIONCONTROL_bus[9];
assign seriesterminationcontrol[10] = sd2a_0_SERIESTERMINATIONCONTROL_bus[10];
assign seriesterminationcontrol[11] = sd2a_0_SERIESTERMINATIONCONTROL_bus[11];
assign seriesterminationcontrol[12] = sd2a_0_SERIESTERMINATIONCONTROL_bus[12];
assign seriesterminationcontrol[13] = sd2a_0_SERIESTERMINATIONCONTROL_bus[13];
assign seriesterminationcontrol[14] = sd2a_0_SERIESTERMINATIONCONTROL_bus[14];
assign seriesterminationcontrol[15] = sd2a_0_SERIESTERMINATIONCONTROL_bus[15];

cyclonev_termination_logic sd2a_0(
	.s2pload(gnd),
	.scanclk(gnd),
	.scanenable(gnd),
	.serdata(\wire_sd1a_serdataout[0] ),
	.enser(4'b0000),
	.parallelterminationcontrol(sd2a_0_PARALLELTERMINATIONCONTROL_bus),
	.seriesterminationcontrol(sd2a_0_SERIESTERMINATIONCONTROL_bus));

cyclonev_termination sd1a_0(
	.clkenusr(gnd),
	.clkusr(gnd),
	.enserusr(gnd),
	.nclrusr(gnd),
	.rzqin(oct_rzqin),
	.scanclk(gnd),
	.scanen(gnd),
	.scanin(gnd),
	.serdatafromcore(gnd),
	.serdatain(gnd),
	.otherenser(10'b0000000000),
	.clkusrdftout(\sd1a_0~O_CLKUSRDFTOUT ),
	.compoutrdn(),
	.compoutrup(),
	.enserout(),
	.scanout(),
	.serdataout(\wire_sd1a_serdataout[0] ),
	.serdatatocore());

endmodule

module Computer_System_hps_sdram_p0 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid_0,
	ctl_reset_n,
	afi_rdata_0,
	afi_rdata_1,
	afi_rdata_2,
	afi_rdata_3,
	afi_rdata_4,
	afi_rdata_5,
	afi_rdata_6,
	afi_rdata_7,
	afi_rdata_8,
	afi_rdata_9,
	afi_rdata_10,
	afi_rdata_11,
	afi_rdata_12,
	afi_rdata_13,
	afi_rdata_14,
	afi_rdata_15,
	afi_rdata_16,
	afi_rdata_17,
	afi_rdata_18,
	afi_rdata_19,
	afi_rdata_20,
	afi_rdata_21,
	afi_rdata_22,
	afi_rdata_23,
	afi_rdata_24,
	afi_rdata_25,
	afi_rdata_26,
	afi_rdata_27,
	afi_rdata_28,
	afi_rdata_29,
	afi_rdata_30,
	afi_rdata_31,
	afi_rdata_32,
	afi_rdata_33,
	afi_rdata_34,
	afi_rdata_35,
	afi_rdata_36,
	afi_rdata_37,
	afi_rdata_38,
	afi_rdata_39,
	afi_rdata_40,
	afi_rdata_41,
	afi_rdata_42,
	afi_rdata_43,
	afi_rdata_44,
	afi_rdata_45,
	afi_rdata_46,
	afi_rdata_47,
	afi_rdata_48,
	afi_rdata_49,
	afi_rdata_50,
	afi_rdata_51,
	afi_rdata_52,
	afi_rdata_53,
	afi_rdata_54,
	afi_rdata_55,
	afi_rdata_56,
	afi_rdata_57,
	afi_rdata_58,
	afi_rdata_59,
	afi_rdata_60,
	afi_rdata_61,
	afi_rdata_62,
	afi_rdata_63,
	afi_rdata_64,
	afi_rdata_65,
	afi_rdata_66,
	afi_rdata_67,
	afi_rdata_68,
	afi_rdata_69,
	afi_rdata_70,
	afi_rdata_71,
	afi_rdata_72,
	afi_rdata_73,
	afi_rdata_74,
	afi_rdata_75,
	afi_rdata_76,
	afi_rdata_77,
	afi_rdata_78,
	afi_rdata_79,
	afi_wlat_0,
	afi_wlat_1,
	afi_wlat_2,
	afi_wlat_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	afi_cas_n_0,
	afi_ras_n_0,
	afi_rst_n_0,
	afi_we_n_0,
	afi_addr_0,
	afi_addr_1,
	afi_addr_2,
	afi_addr_3,
	afi_addr_4,
	afi_addr_5,
	afi_addr_6,
	afi_addr_7,
	afi_addr_8,
	afi_addr_9,
	afi_addr_10,
	afi_addr_11,
	afi_addr_12,
	afi_addr_13,
	afi_addr_14,
	afi_addr_15,
	afi_addr_16,
	afi_addr_17,
	afi_addr_18,
	afi_addr_19,
	afi_ba_0,
	afi_ba_1,
	afi_ba_2,
	afi_cke_0,
	afi_cke_1,
	afi_cs_n_0,
	afi_cs_n_1,
	afi_dm_int_0,
	afi_dm_int_1,
	afi_dm_int_2,
	afi_dm_int_3,
	afi_dm_int_4,
	afi_dm_int_5,
	afi_dm_int_6,
	afi_dm_int_7,
	afi_dm_int_8,
	afi_dm_int_9,
	afi_dqs_burst_0,
	afi_dqs_burst_1,
	afi_dqs_burst_2,
	afi_dqs_burst_3,
	afi_dqs_burst_4,
	afi_odt_0,
	afi_odt_1,
	afi_rdata_en_0,
	afi_rdata_en_1,
	afi_rdata_en_2,
	afi_rdata_en_3,
	afi_rdata_en_4,
	afi_rdata_en_full_0,
	afi_rdata_en_full_1,
	afi_rdata_en_full_2,
	afi_rdata_en_full_3,
	afi_rdata_en_full_4,
	afi_wdata_int_0,
	afi_wdata_int_1,
	afi_wdata_int_2,
	afi_wdata_int_3,
	afi_wdata_int_4,
	afi_wdata_int_5,
	afi_wdata_int_6,
	afi_wdata_int_7,
	afi_wdata_int_8,
	afi_wdata_int_9,
	afi_wdata_int_10,
	afi_wdata_int_11,
	afi_wdata_int_12,
	afi_wdata_int_13,
	afi_wdata_int_14,
	afi_wdata_int_15,
	afi_wdata_int_16,
	afi_wdata_int_17,
	afi_wdata_int_18,
	afi_wdata_int_19,
	afi_wdata_int_20,
	afi_wdata_int_21,
	afi_wdata_int_22,
	afi_wdata_int_23,
	afi_wdata_int_24,
	afi_wdata_int_25,
	afi_wdata_int_26,
	afi_wdata_int_27,
	afi_wdata_int_28,
	afi_wdata_int_29,
	afi_wdata_int_30,
	afi_wdata_int_31,
	afi_wdata_int_32,
	afi_wdata_int_33,
	afi_wdata_int_34,
	afi_wdata_int_35,
	afi_wdata_int_36,
	afi_wdata_int_37,
	afi_wdata_int_38,
	afi_wdata_int_39,
	afi_wdata_int_40,
	afi_wdata_int_41,
	afi_wdata_int_42,
	afi_wdata_int_43,
	afi_wdata_int_44,
	afi_wdata_int_45,
	afi_wdata_int_46,
	afi_wdata_int_47,
	afi_wdata_int_48,
	afi_wdata_int_49,
	afi_wdata_int_50,
	afi_wdata_int_51,
	afi_wdata_int_52,
	afi_wdata_int_53,
	afi_wdata_int_54,
	afi_wdata_int_55,
	afi_wdata_int_56,
	afi_wdata_int_57,
	afi_wdata_int_58,
	afi_wdata_int_59,
	afi_wdata_int_60,
	afi_wdata_int_61,
	afi_wdata_int_62,
	afi_wdata_int_63,
	afi_wdata_int_64,
	afi_wdata_int_65,
	afi_wdata_int_66,
	afi_wdata_int_67,
	afi_wdata_int_68,
	afi_wdata_int_69,
	afi_wdata_int_70,
	afi_wdata_int_71,
	afi_wdata_int_72,
	afi_wdata_int_73,
	afi_wdata_int_74,
	afi_wdata_int_75,
	afi_wdata_int_76,
	afi_wdata_int_77,
	afi_wdata_int_78,
	afi_wdata_int_79,
	afi_wdata_valid_0,
	afi_wdata_valid_1,
	afi_wdata_valid_2,
	afi_wdata_valid_3,
	afi_wdata_valid_4,
	cfg_addlat_wire_0,
	cfg_addlat_wire_1,
	cfg_addlat_wire_2,
	cfg_addlat_wire_3,
	cfg_addlat_wire_4,
	cfg_bankaddrwidth_wire_0,
	cfg_bankaddrwidth_wire_1,
	cfg_bankaddrwidth_wire_2,
	cfg_caswrlat_wire_0,
	cfg_caswrlat_wire_1,
	cfg_caswrlat_wire_2,
	cfg_caswrlat_wire_3,
	cfg_coladdrwidth_wire_0,
	cfg_coladdrwidth_wire_1,
	cfg_coladdrwidth_wire_2,
	cfg_coladdrwidth_wire_3,
	cfg_coladdrwidth_wire_4,
	cfg_csaddrwidth_wire_0,
	cfg_csaddrwidth_wire_1,
	cfg_csaddrwidth_wire_2,
	cfg_devicewidth_wire_0,
	cfg_devicewidth_wire_1,
	cfg_devicewidth_wire_2,
	cfg_devicewidth_wire_3,
	cfg_interfacewidth_wire_0,
	cfg_interfacewidth_wire_1,
	cfg_interfacewidth_wire_2,
	cfg_interfacewidth_wire_3,
	cfg_interfacewidth_wire_4,
	cfg_interfacewidth_wire_5,
	cfg_interfacewidth_wire_6,
	cfg_interfacewidth_wire_7,
	cfg_rowaddrwidth_wire_0,
	cfg_rowaddrwidth_wire_1,
	cfg_rowaddrwidth_wire_2,
	cfg_rowaddrwidth_wire_3,
	cfg_rowaddrwidth_wire_4,
	cfg_tcl_wire_0,
	cfg_tcl_wire_1,
	cfg_tcl_wire_2,
	cfg_tcl_wire_3,
	cfg_tcl_wire_4,
	cfg_tmrd_wire_0,
	cfg_tmrd_wire_1,
	cfg_tmrd_wire_2,
	cfg_tmrd_wire_3,
	cfg_trefi_wire_0,
	cfg_trefi_wire_1,
	cfg_trefi_wire_2,
	cfg_trefi_wire_3,
	cfg_trefi_wire_4,
	cfg_trefi_wire_5,
	cfg_trefi_wire_6,
	cfg_trefi_wire_7,
	cfg_trefi_wire_8,
	cfg_trefi_wire_9,
	cfg_trefi_wire_10,
	cfg_trefi_wire_11,
	cfg_trefi_wire_12,
	cfg_trfc_wire_0,
	cfg_trfc_wire_1,
	cfg_trfc_wire_2,
	cfg_trfc_wire_3,
	cfg_trfc_wire_4,
	cfg_trfc_wire_5,
	cfg_trfc_wire_6,
	cfg_trfc_wire_7,
	cfg_twr_wire_0,
	cfg_twr_wire_1,
	cfg_twr_wire_2,
	cfg_twr_wire_3,
	afi_mem_clk_disable_0,
	cfg_dramconfig_wire_0,
	cfg_dramconfig_wire_1,
	cfg_dramconfig_wire_2,
	cfg_dramconfig_wire_3,
	cfg_dramconfig_wire_4,
	cfg_dramconfig_wire_5,
	cfg_dramconfig_wire_6,
	cfg_dramconfig_wire_7,
	cfg_dramconfig_wire_8,
	cfg_dramconfig_wire_9,
	cfg_dramconfig_wire_10,
	cfg_dramconfig_wire_11,
	cfg_dramconfig_wire_12,
	cfg_dramconfig_wire_13,
	cfg_dramconfig_wire_14,
	cfg_dramconfig_wire_15,
	cfg_dramconfig_wire_16,
	cfg_dramconfig_wire_17,
	cfg_dramconfig_wire_18,
	cfg_dramconfig_wire_19,
	cfg_dramconfig_wire_20,
	ctl_clk,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	afi_cal_fail;
output 	afi_cal_success;
output 	afi_rdata_valid_0;
output 	ctl_reset_n;
output 	afi_rdata_0;
output 	afi_rdata_1;
output 	afi_rdata_2;
output 	afi_rdata_3;
output 	afi_rdata_4;
output 	afi_rdata_5;
output 	afi_rdata_6;
output 	afi_rdata_7;
output 	afi_rdata_8;
output 	afi_rdata_9;
output 	afi_rdata_10;
output 	afi_rdata_11;
output 	afi_rdata_12;
output 	afi_rdata_13;
output 	afi_rdata_14;
output 	afi_rdata_15;
output 	afi_rdata_16;
output 	afi_rdata_17;
output 	afi_rdata_18;
output 	afi_rdata_19;
output 	afi_rdata_20;
output 	afi_rdata_21;
output 	afi_rdata_22;
output 	afi_rdata_23;
output 	afi_rdata_24;
output 	afi_rdata_25;
output 	afi_rdata_26;
output 	afi_rdata_27;
output 	afi_rdata_28;
output 	afi_rdata_29;
output 	afi_rdata_30;
output 	afi_rdata_31;
output 	afi_rdata_32;
output 	afi_rdata_33;
output 	afi_rdata_34;
output 	afi_rdata_35;
output 	afi_rdata_36;
output 	afi_rdata_37;
output 	afi_rdata_38;
output 	afi_rdata_39;
output 	afi_rdata_40;
output 	afi_rdata_41;
output 	afi_rdata_42;
output 	afi_rdata_43;
output 	afi_rdata_44;
output 	afi_rdata_45;
output 	afi_rdata_46;
output 	afi_rdata_47;
output 	afi_rdata_48;
output 	afi_rdata_49;
output 	afi_rdata_50;
output 	afi_rdata_51;
output 	afi_rdata_52;
output 	afi_rdata_53;
output 	afi_rdata_54;
output 	afi_rdata_55;
output 	afi_rdata_56;
output 	afi_rdata_57;
output 	afi_rdata_58;
output 	afi_rdata_59;
output 	afi_rdata_60;
output 	afi_rdata_61;
output 	afi_rdata_62;
output 	afi_rdata_63;
output 	afi_rdata_64;
output 	afi_rdata_65;
output 	afi_rdata_66;
output 	afi_rdata_67;
output 	afi_rdata_68;
output 	afi_rdata_69;
output 	afi_rdata_70;
output 	afi_rdata_71;
output 	afi_rdata_72;
output 	afi_rdata_73;
output 	afi_rdata_74;
output 	afi_rdata_75;
output 	afi_rdata_76;
output 	afi_rdata_77;
output 	afi_rdata_78;
output 	afi_rdata_79;
output 	afi_wlat_0;
output 	afi_wlat_1;
output 	afi_wlat_2;
output 	afi_wlat_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	afi_cas_n_0;
input 	afi_ras_n_0;
input 	afi_rst_n_0;
input 	afi_we_n_0;
input 	afi_addr_0;
input 	afi_addr_1;
input 	afi_addr_2;
input 	afi_addr_3;
input 	afi_addr_4;
input 	afi_addr_5;
input 	afi_addr_6;
input 	afi_addr_7;
input 	afi_addr_8;
input 	afi_addr_9;
input 	afi_addr_10;
input 	afi_addr_11;
input 	afi_addr_12;
input 	afi_addr_13;
input 	afi_addr_14;
input 	afi_addr_15;
input 	afi_addr_16;
input 	afi_addr_17;
input 	afi_addr_18;
input 	afi_addr_19;
input 	afi_ba_0;
input 	afi_ba_1;
input 	afi_ba_2;
input 	afi_cke_0;
input 	afi_cke_1;
input 	afi_cs_n_0;
input 	afi_cs_n_1;
input 	afi_dm_int_0;
input 	afi_dm_int_1;
input 	afi_dm_int_2;
input 	afi_dm_int_3;
input 	afi_dm_int_4;
input 	afi_dm_int_5;
input 	afi_dm_int_6;
input 	afi_dm_int_7;
input 	afi_dm_int_8;
input 	afi_dm_int_9;
input 	afi_dqs_burst_0;
input 	afi_dqs_burst_1;
input 	afi_dqs_burst_2;
input 	afi_dqs_burst_3;
input 	afi_dqs_burst_4;
input 	afi_odt_0;
input 	afi_odt_1;
input 	afi_rdata_en_0;
input 	afi_rdata_en_1;
input 	afi_rdata_en_2;
input 	afi_rdata_en_3;
input 	afi_rdata_en_4;
input 	afi_rdata_en_full_0;
input 	afi_rdata_en_full_1;
input 	afi_rdata_en_full_2;
input 	afi_rdata_en_full_3;
input 	afi_rdata_en_full_4;
input 	afi_wdata_int_0;
input 	afi_wdata_int_1;
input 	afi_wdata_int_2;
input 	afi_wdata_int_3;
input 	afi_wdata_int_4;
input 	afi_wdata_int_5;
input 	afi_wdata_int_6;
input 	afi_wdata_int_7;
input 	afi_wdata_int_8;
input 	afi_wdata_int_9;
input 	afi_wdata_int_10;
input 	afi_wdata_int_11;
input 	afi_wdata_int_12;
input 	afi_wdata_int_13;
input 	afi_wdata_int_14;
input 	afi_wdata_int_15;
input 	afi_wdata_int_16;
input 	afi_wdata_int_17;
input 	afi_wdata_int_18;
input 	afi_wdata_int_19;
input 	afi_wdata_int_20;
input 	afi_wdata_int_21;
input 	afi_wdata_int_22;
input 	afi_wdata_int_23;
input 	afi_wdata_int_24;
input 	afi_wdata_int_25;
input 	afi_wdata_int_26;
input 	afi_wdata_int_27;
input 	afi_wdata_int_28;
input 	afi_wdata_int_29;
input 	afi_wdata_int_30;
input 	afi_wdata_int_31;
input 	afi_wdata_int_32;
input 	afi_wdata_int_33;
input 	afi_wdata_int_34;
input 	afi_wdata_int_35;
input 	afi_wdata_int_36;
input 	afi_wdata_int_37;
input 	afi_wdata_int_38;
input 	afi_wdata_int_39;
input 	afi_wdata_int_40;
input 	afi_wdata_int_41;
input 	afi_wdata_int_42;
input 	afi_wdata_int_43;
input 	afi_wdata_int_44;
input 	afi_wdata_int_45;
input 	afi_wdata_int_46;
input 	afi_wdata_int_47;
input 	afi_wdata_int_48;
input 	afi_wdata_int_49;
input 	afi_wdata_int_50;
input 	afi_wdata_int_51;
input 	afi_wdata_int_52;
input 	afi_wdata_int_53;
input 	afi_wdata_int_54;
input 	afi_wdata_int_55;
input 	afi_wdata_int_56;
input 	afi_wdata_int_57;
input 	afi_wdata_int_58;
input 	afi_wdata_int_59;
input 	afi_wdata_int_60;
input 	afi_wdata_int_61;
input 	afi_wdata_int_62;
input 	afi_wdata_int_63;
input 	afi_wdata_int_64;
input 	afi_wdata_int_65;
input 	afi_wdata_int_66;
input 	afi_wdata_int_67;
input 	afi_wdata_int_68;
input 	afi_wdata_int_69;
input 	afi_wdata_int_70;
input 	afi_wdata_int_71;
input 	afi_wdata_int_72;
input 	afi_wdata_int_73;
input 	afi_wdata_int_74;
input 	afi_wdata_int_75;
input 	afi_wdata_int_76;
input 	afi_wdata_int_77;
input 	afi_wdata_int_78;
input 	afi_wdata_int_79;
input 	afi_wdata_valid_0;
input 	afi_wdata_valid_1;
input 	afi_wdata_valid_2;
input 	afi_wdata_valid_3;
input 	afi_wdata_valid_4;
input 	cfg_addlat_wire_0;
input 	cfg_addlat_wire_1;
input 	cfg_addlat_wire_2;
input 	cfg_addlat_wire_3;
input 	cfg_addlat_wire_4;
input 	cfg_bankaddrwidth_wire_0;
input 	cfg_bankaddrwidth_wire_1;
input 	cfg_bankaddrwidth_wire_2;
input 	cfg_caswrlat_wire_0;
input 	cfg_caswrlat_wire_1;
input 	cfg_caswrlat_wire_2;
input 	cfg_caswrlat_wire_3;
input 	cfg_coladdrwidth_wire_0;
input 	cfg_coladdrwidth_wire_1;
input 	cfg_coladdrwidth_wire_2;
input 	cfg_coladdrwidth_wire_3;
input 	cfg_coladdrwidth_wire_4;
input 	cfg_csaddrwidth_wire_0;
input 	cfg_csaddrwidth_wire_1;
input 	cfg_csaddrwidth_wire_2;
input 	cfg_devicewidth_wire_0;
input 	cfg_devicewidth_wire_1;
input 	cfg_devicewidth_wire_2;
input 	cfg_devicewidth_wire_3;
input 	cfg_interfacewidth_wire_0;
input 	cfg_interfacewidth_wire_1;
input 	cfg_interfacewidth_wire_2;
input 	cfg_interfacewidth_wire_3;
input 	cfg_interfacewidth_wire_4;
input 	cfg_interfacewidth_wire_5;
input 	cfg_interfacewidth_wire_6;
input 	cfg_interfacewidth_wire_7;
input 	cfg_rowaddrwidth_wire_0;
input 	cfg_rowaddrwidth_wire_1;
input 	cfg_rowaddrwidth_wire_2;
input 	cfg_rowaddrwidth_wire_3;
input 	cfg_rowaddrwidth_wire_4;
input 	cfg_tcl_wire_0;
input 	cfg_tcl_wire_1;
input 	cfg_tcl_wire_2;
input 	cfg_tcl_wire_3;
input 	cfg_tcl_wire_4;
input 	cfg_tmrd_wire_0;
input 	cfg_tmrd_wire_1;
input 	cfg_tmrd_wire_2;
input 	cfg_tmrd_wire_3;
input 	cfg_trefi_wire_0;
input 	cfg_trefi_wire_1;
input 	cfg_trefi_wire_2;
input 	cfg_trefi_wire_3;
input 	cfg_trefi_wire_4;
input 	cfg_trefi_wire_5;
input 	cfg_trefi_wire_6;
input 	cfg_trefi_wire_7;
input 	cfg_trefi_wire_8;
input 	cfg_trefi_wire_9;
input 	cfg_trefi_wire_10;
input 	cfg_trefi_wire_11;
input 	cfg_trefi_wire_12;
input 	cfg_trfc_wire_0;
input 	cfg_trfc_wire_1;
input 	cfg_trfc_wire_2;
input 	cfg_trfc_wire_3;
input 	cfg_trfc_wire_4;
input 	cfg_trfc_wire_5;
input 	cfg_trfc_wire_6;
input 	cfg_trfc_wire_7;
input 	cfg_twr_wire_0;
input 	cfg_twr_wire_1;
input 	cfg_twr_wire_2;
input 	cfg_twr_wire_3;
input 	afi_mem_clk_disable_0;
input 	cfg_dramconfig_wire_0;
input 	cfg_dramconfig_wire_1;
input 	cfg_dramconfig_wire_2;
input 	cfg_dramconfig_wire_3;
input 	cfg_dramconfig_wire_4;
input 	cfg_dramconfig_wire_5;
input 	cfg_dramconfig_wire_6;
input 	cfg_dramconfig_wire_7;
input 	cfg_dramconfig_wire_8;
input 	cfg_dramconfig_wire_9;
input 	cfg_dramconfig_wire_10;
input 	cfg_dramconfig_wire_11;
input 	cfg_dramconfig_wire_12;
input 	cfg_dramconfig_wire_13;
input 	cfg_dramconfig_wire_14;
input 	cfg_dramconfig_wire_15;
input 	cfg_dramconfig_wire_16;
input 	cfg_dramconfig_wire_17;
input 	cfg_dramconfig_wire_18;
input 	cfg_dramconfig_wire_19;
input 	cfg_dramconfig_wire_20;
output 	ctl_clk;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_hps_sdram_p0_acv_hard_memphy umemphy(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.afi_cal_fail(afi_cal_fail),
	.afi_cal_success(afi_cal_success),
	.afi_rdata_valid({afi_rdata_valid_0}),
	.ctl_reset_n(ctl_reset_n),
	.afi_rdata({afi_rdata_79,afi_rdata_78,afi_rdata_77,afi_rdata_76,afi_rdata_75,afi_rdata_74,afi_rdata_73,afi_rdata_72,afi_rdata_71,afi_rdata_70,afi_rdata_69,afi_rdata_68,afi_rdata_67,afi_rdata_66,afi_rdata_65,afi_rdata_64,afi_rdata_63,afi_rdata_62,afi_rdata_61,afi_rdata_60,afi_rdata_59,
afi_rdata_58,afi_rdata_57,afi_rdata_56,afi_rdata_55,afi_rdata_54,afi_rdata_53,afi_rdata_52,afi_rdata_51,afi_rdata_50,afi_rdata_49,afi_rdata_48,afi_rdata_47,afi_rdata_46,afi_rdata_45,afi_rdata_44,afi_rdata_43,afi_rdata_42,afi_rdata_41,afi_rdata_40,afi_rdata_39,afi_rdata_38,
afi_rdata_37,afi_rdata_36,afi_rdata_35,afi_rdata_34,afi_rdata_33,afi_rdata_32,afi_rdata_31,afi_rdata_30,afi_rdata_29,afi_rdata_28,afi_rdata_27,afi_rdata_26,afi_rdata_25,afi_rdata_24,afi_rdata_23,afi_rdata_22,afi_rdata_21,afi_rdata_20,afi_rdata_19,afi_rdata_18,afi_rdata_17,
afi_rdata_16,afi_rdata_15,afi_rdata_14,afi_rdata_13,afi_rdata_12,afi_rdata_11,afi_rdata_10,afi_rdata_9,afi_rdata_8,afi_rdata_7,afi_rdata_6,afi_rdata_5,afi_rdata_4,afi_rdata_3,afi_rdata_2,afi_rdata_1,afi_rdata_0}),
	.afi_wlat({afi_wlat_3,afi_wlat_2,afi_wlat_1,afi_wlat_0}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.afi_cas_n({afi_cas_n_0}),
	.afi_ras_n({afi_ras_n_0}),
	.afi_rst_n({afi_rst_n_0}),
	.afi_we_n({afi_we_n_0}),
	.afi_addr({afi_addr_19,afi_addr_18,afi_addr_17,afi_addr_16,afi_addr_15,afi_addr_14,afi_addr_13,afi_addr_12,afi_addr_11,afi_addr_10,afi_addr_9,afi_addr_8,afi_addr_7,afi_addr_6,afi_addr_5,afi_addr_4,afi_addr_3,afi_addr_2,afi_addr_1,afi_addr_0}),
	.afi_ba({afi_ba_2,afi_ba_1,afi_ba_0}),
	.afi_cke({afi_cke_1,afi_cke_0}),
	.afi_cs_n({afi_cs_n_1,afi_cs_n_0}),
	.afi_dm({afi_dm_int_9,afi_dm_int_8,afi_dm_int_7,afi_dm_int_6,afi_dm_int_5,afi_dm_int_4,afi_dm_int_3,afi_dm_int_2,afi_dm_int_1,afi_dm_int_0}),
	.afi_dqs_burst({afi_dqs_burst_4,afi_dqs_burst_3,afi_dqs_burst_2,afi_dqs_burst_1,afi_dqs_burst_0}),
	.afi_odt({afi_odt_1,afi_odt_0}),
	.afi_rdata_en({afi_rdata_en_4,afi_rdata_en_3,afi_rdata_en_2,afi_rdata_en_1,afi_rdata_en_0}),
	.afi_rdata_en_full({afi_rdata_en_full_4,afi_rdata_en_full_3,afi_rdata_en_full_2,afi_rdata_en_full_1,afi_rdata_en_full_0}),
	.afi_wdata({afi_wdata_int_79,afi_wdata_int_78,afi_wdata_int_77,afi_wdata_int_76,afi_wdata_int_75,afi_wdata_int_74,afi_wdata_int_73,afi_wdata_int_72,afi_wdata_int_71,afi_wdata_int_70,afi_wdata_int_69,afi_wdata_int_68,afi_wdata_int_67,afi_wdata_int_66,afi_wdata_int_65,afi_wdata_int_64,
afi_wdata_int_63,afi_wdata_int_62,afi_wdata_int_61,afi_wdata_int_60,afi_wdata_int_59,afi_wdata_int_58,afi_wdata_int_57,afi_wdata_int_56,afi_wdata_int_55,afi_wdata_int_54,afi_wdata_int_53,afi_wdata_int_52,afi_wdata_int_51,afi_wdata_int_50,afi_wdata_int_49,afi_wdata_int_48,
afi_wdata_int_47,afi_wdata_int_46,afi_wdata_int_45,afi_wdata_int_44,afi_wdata_int_43,afi_wdata_int_42,afi_wdata_int_41,afi_wdata_int_40,afi_wdata_int_39,afi_wdata_int_38,afi_wdata_int_37,afi_wdata_int_36,afi_wdata_int_35,afi_wdata_int_34,afi_wdata_int_33,afi_wdata_int_32,
afi_wdata_int_31,afi_wdata_int_30,afi_wdata_int_29,afi_wdata_int_28,afi_wdata_int_27,afi_wdata_int_26,afi_wdata_int_25,afi_wdata_int_24,afi_wdata_int_23,afi_wdata_int_22,afi_wdata_int_21,afi_wdata_int_20,afi_wdata_int_19,afi_wdata_int_18,afi_wdata_int_17,afi_wdata_int_16,
afi_wdata_int_15,afi_wdata_int_14,afi_wdata_int_13,afi_wdata_int_12,afi_wdata_int_11,afi_wdata_int_10,afi_wdata_int_9,afi_wdata_int_8,afi_wdata_int_7,afi_wdata_int_6,afi_wdata_int_5,afi_wdata_int_4,afi_wdata_int_3,afi_wdata_int_2,afi_wdata_int_1,afi_wdata_int_0}),
	.afi_wdata_valid({afi_wdata_valid_4,afi_wdata_valid_3,afi_wdata_valid_2,afi_wdata_valid_1,afi_wdata_valid_0}),
	.cfg_addlat({gnd,gnd,gnd,cfg_addlat_wire_4,cfg_addlat_wire_3,cfg_addlat_wire_2,cfg_addlat_wire_1,cfg_addlat_wire_0}),
	.cfg_bankaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_bankaddrwidth_wire_2,cfg_bankaddrwidth_wire_1,cfg_bankaddrwidth_wire_0}),
	.cfg_caswrlat({gnd,gnd,gnd,gnd,cfg_caswrlat_wire_3,cfg_caswrlat_wire_2,cfg_caswrlat_wire_1,cfg_caswrlat_wire_0}),
	.cfg_coladdrwidth({gnd,gnd,gnd,cfg_coladdrwidth_wire_4,cfg_coladdrwidth_wire_3,cfg_coladdrwidth_wire_2,cfg_coladdrwidth_wire_1,cfg_coladdrwidth_wire_0}),
	.cfg_csaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_csaddrwidth_wire_2,cfg_csaddrwidth_wire_1,cfg_csaddrwidth_wire_0}),
	.cfg_devicewidth({gnd,gnd,gnd,gnd,cfg_devicewidth_wire_3,cfg_devicewidth_wire_2,cfg_devicewidth_wire_1,cfg_devicewidth_wire_0}),
	.cfg_interfacewidth({cfg_interfacewidth_wire_7,cfg_interfacewidth_wire_6,cfg_interfacewidth_wire_5,cfg_interfacewidth_wire_4,cfg_interfacewidth_wire_3,cfg_interfacewidth_wire_2,cfg_interfacewidth_wire_1,cfg_interfacewidth_wire_0}),
	.cfg_rowaddrwidth({gnd,gnd,gnd,cfg_rowaddrwidth_wire_4,cfg_rowaddrwidth_wire_3,cfg_rowaddrwidth_wire_2,cfg_rowaddrwidth_wire_1,cfg_rowaddrwidth_wire_0}),
	.cfg_tcl({gnd,gnd,gnd,cfg_tcl_wire_4,cfg_tcl_wire_3,cfg_tcl_wire_2,cfg_tcl_wire_1,cfg_tcl_wire_0}),
	.cfg_tmrd({gnd,gnd,gnd,gnd,cfg_tmrd_wire_3,cfg_tmrd_wire_2,cfg_tmrd_wire_1,cfg_tmrd_wire_0}),
	.cfg_trefi({gnd,gnd,gnd,cfg_trefi_wire_12,cfg_trefi_wire_11,cfg_trefi_wire_10,cfg_trefi_wire_9,cfg_trefi_wire_8,cfg_trefi_wire_7,cfg_trefi_wire_6,cfg_trefi_wire_5,cfg_trefi_wire_4,cfg_trefi_wire_3,cfg_trefi_wire_2,cfg_trefi_wire_1,cfg_trefi_wire_0}),
	.cfg_trfc({cfg_trfc_wire_7,cfg_trfc_wire_6,cfg_trfc_wire_5,cfg_trfc_wire_4,cfg_trfc_wire_3,cfg_trfc_wire_2,cfg_trfc_wire_1,cfg_trfc_wire_0}),
	.cfg_twr({gnd,gnd,gnd,gnd,cfg_twr_wire_3,cfg_twr_wire_2,cfg_twr_wire_1,cfg_twr_wire_0}),
	.afi_mem_clk_disable({afi_mem_clk_disable_0}),
	.cfg_dramconfig({gnd,gnd,gnd,cfg_dramconfig_wire_20,cfg_dramconfig_wire_19,cfg_dramconfig_wire_18,cfg_dramconfig_wire_17,cfg_dramconfig_wire_16,cfg_dramconfig_wire_15,cfg_dramconfig_wire_14,cfg_dramconfig_wire_13,cfg_dramconfig_wire_12,cfg_dramconfig_wire_11,cfg_dramconfig_wire_10,
cfg_dramconfig_wire_9,cfg_dramconfig_wire_8,cfg_dramconfig_wire_7,cfg_dramconfig_wire_6,cfg_dramconfig_wire_5,cfg_dramconfig_wire_4,cfg_dramconfig_wire_3,cfg_dramconfig_wire_2,cfg_dramconfig_wire_1,cfg_dramconfig_wire_0}),
	.ctl_clk(ctl_clk),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

endmodule

module Computer_System_hps_sdram_p0_acv_hard_memphy (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid,
	ctl_reset_n,
	afi_rdata,
	afi_wlat,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	afi_cas_n,
	afi_ras_n,
	afi_rst_n,
	afi_we_n,
	afi_addr,
	afi_ba,
	afi_cke,
	afi_cs_n,
	afi_dm,
	afi_dqs_burst,
	afi_odt,
	afi_rdata_en,
	afi_rdata_en_full,
	afi_wdata,
	afi_wdata_valid,
	cfg_addlat,
	cfg_bankaddrwidth,
	cfg_caswrlat,
	cfg_coladdrwidth,
	cfg_csaddrwidth,
	cfg_devicewidth,
	cfg_interfacewidth,
	cfg_rowaddrwidth,
	cfg_tcl,
	cfg_tmrd,
	cfg_trefi,
	cfg_trfc,
	cfg_twr,
	afi_mem_clk_disable,
	cfg_dramconfig,
	ctl_clk,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	afi_cal_fail;
output 	afi_cal_success;
output 	[0:0] afi_rdata_valid;
output 	ctl_reset_n;
output 	[79:0] afi_rdata;
output 	[3:0] afi_wlat;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	[0:0] afi_cas_n;
input 	[0:0] afi_ras_n;
input 	[0:0] afi_rst_n;
input 	[0:0] afi_we_n;
input 	[19:0] afi_addr;
input 	[2:0] afi_ba;
input 	[1:0] afi_cke;
input 	[1:0] afi_cs_n;
input 	[9:0] afi_dm;
input 	[4:0] afi_dqs_burst;
input 	[1:0] afi_odt;
input 	[4:0] afi_rdata_en;
input 	[4:0] afi_rdata_en_full;
input 	[79:0] afi_wdata;
input 	[4:0] afi_wdata_valid;
input 	[7:0] cfg_addlat;
input 	[7:0] cfg_bankaddrwidth;
input 	[7:0] cfg_caswrlat;
input 	[7:0] cfg_coladdrwidth;
input 	[7:0] cfg_csaddrwidth;
input 	[7:0] cfg_devicewidth;
input 	[7:0] cfg_interfacewidth;
input 	[7:0] cfg_rowaddrwidth;
input 	[7:0] cfg_tcl;
input 	[7:0] cfg_tmrd;
input 	[15:0] cfg_trefi;
input 	[7:0] cfg_trfc;
input 	[7:0] cfg_twr;
input 	[0:0] afi_mem_clk_disable;
input 	[23:0] cfg_dramconfig;
output 	ctl_clk;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \memphy_ldc|leveled_hr_clocks[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \phy_ddio_address[0] ;
wire \phy_ddio_address[1] ;
wire \phy_ddio_address[2] ;
wire \phy_ddio_address[3] ;
wire \phy_ddio_address[4] ;
wire \phy_ddio_address[5] ;
wire \phy_ddio_address[6] ;
wire \phy_ddio_address[7] ;
wire \phy_ddio_address[8] ;
wire \phy_ddio_address[9] ;
wire \phy_ddio_address[10] ;
wire \phy_ddio_address[11] ;
wire \phy_ddio_address[12] ;
wire \phy_ddio_address[13] ;
wire \phy_ddio_address[14] ;
wire \phy_ddio_address[15] ;
wire \phy_ddio_address[16] ;
wire \phy_ddio_address[17] ;
wire \phy_ddio_address[18] ;
wire \phy_ddio_address[19] ;
wire \phy_ddio_address[20] ;
wire \phy_ddio_address[21] ;
wire \phy_ddio_address[22] ;
wire \phy_ddio_address[23] ;
wire \phy_ddio_address[24] ;
wire \phy_ddio_address[25] ;
wire \phy_ddio_address[26] ;
wire \phy_ddio_address[27] ;
wire \phy_ddio_address[28] ;
wire \phy_ddio_address[29] ;
wire \phy_ddio_address[30] ;
wire \phy_ddio_address[31] ;
wire \phy_ddio_address[32] ;
wire \phy_ddio_address[33] ;
wire \phy_ddio_address[34] ;
wire \phy_ddio_address[35] ;
wire \phy_ddio_address[36] ;
wire \phy_ddio_address[37] ;
wire \phy_ddio_address[38] ;
wire \phy_ddio_address[39] ;
wire \phy_ddio_address[40] ;
wire \phy_ddio_address[41] ;
wire \phy_ddio_address[42] ;
wire \phy_ddio_address[43] ;
wire \phy_ddio_address[44] ;
wire \phy_ddio_address[45] ;
wire \phy_ddio_address[46] ;
wire \phy_ddio_address[47] ;
wire \phy_ddio_address[48] ;
wire \phy_ddio_address[49] ;
wire \phy_ddio_address[50] ;
wire \phy_ddio_address[51] ;
wire \phy_ddio_address[52] ;
wire \phy_ddio_address[53] ;
wire \phy_ddio_address[54] ;
wire \phy_ddio_address[55] ;
wire \phy_ddio_address[56] ;
wire \phy_ddio_address[57] ;
wire \phy_ddio_address[58] ;
wire \phy_ddio_address[59] ;
wire \phy_ddio_bank[0] ;
wire \phy_ddio_bank[1] ;
wire \phy_ddio_bank[2] ;
wire \phy_ddio_bank[3] ;
wire \phy_ddio_bank[4] ;
wire \phy_ddio_bank[5] ;
wire \phy_ddio_bank[6] ;
wire \phy_ddio_bank[7] ;
wire \phy_ddio_bank[8] ;
wire \phy_ddio_bank[9] ;
wire \phy_ddio_bank[10] ;
wire \phy_ddio_bank[11] ;
wire \phy_ddio_cas_n[0] ;
wire \phy_ddio_cas_n[1] ;
wire \phy_ddio_cas_n[2] ;
wire \phy_ddio_cas_n[3] ;
wire \phy_ddio_ck[0] ;
wire \phy_ddio_ck[1] ;
wire \phy_ddio_cke[0] ;
wire \phy_ddio_cke[1] ;
wire \phy_ddio_cke[2] ;
wire \phy_ddio_cke[3] ;
wire \phy_ddio_cs_n[0] ;
wire \phy_ddio_cs_n[1] ;
wire \phy_ddio_cs_n[2] ;
wire \phy_ddio_cs_n[3] ;
wire \phy_ddio_dmdout[0] ;
wire \phy_ddio_dmdout[1] ;
wire \phy_ddio_dmdout[2] ;
wire \phy_ddio_dmdout[3] ;
wire \phy_ddio_dmdout[4] ;
wire \phy_ddio_dmdout[5] ;
wire \phy_ddio_dmdout[6] ;
wire \phy_ddio_dmdout[7] ;
wire \phy_ddio_dmdout[8] ;
wire \phy_ddio_dmdout[9] ;
wire \phy_ddio_dmdout[10] ;
wire \phy_ddio_dmdout[11] ;
wire \phy_ddio_dmdout[12] ;
wire \phy_ddio_dmdout[13] ;
wire \phy_ddio_dmdout[14] ;
wire \phy_ddio_dmdout[15] ;
wire \phy_ddio_dqdout[0] ;
wire \phy_ddio_dqdout[1] ;
wire \phy_ddio_dqdout[2] ;
wire \phy_ddio_dqdout[3] ;
wire \phy_ddio_dqdout[4] ;
wire \phy_ddio_dqdout[5] ;
wire \phy_ddio_dqdout[6] ;
wire \phy_ddio_dqdout[7] ;
wire \phy_ddio_dqdout[8] ;
wire \phy_ddio_dqdout[9] ;
wire \phy_ddio_dqdout[10] ;
wire \phy_ddio_dqdout[11] ;
wire \phy_ddio_dqdout[12] ;
wire \phy_ddio_dqdout[13] ;
wire \phy_ddio_dqdout[14] ;
wire \phy_ddio_dqdout[15] ;
wire \phy_ddio_dqdout[16] ;
wire \phy_ddio_dqdout[17] ;
wire \phy_ddio_dqdout[18] ;
wire \phy_ddio_dqdout[19] ;
wire \phy_ddio_dqdout[20] ;
wire \phy_ddio_dqdout[21] ;
wire \phy_ddio_dqdout[22] ;
wire \phy_ddio_dqdout[23] ;
wire \phy_ddio_dqdout[24] ;
wire \phy_ddio_dqdout[25] ;
wire \phy_ddio_dqdout[26] ;
wire \phy_ddio_dqdout[27] ;
wire \phy_ddio_dqdout[28] ;
wire \phy_ddio_dqdout[29] ;
wire \phy_ddio_dqdout[30] ;
wire \phy_ddio_dqdout[31] ;
wire \phy_ddio_dqdout[36] ;
wire \phy_ddio_dqdout[37] ;
wire \phy_ddio_dqdout[38] ;
wire \phy_ddio_dqdout[39] ;
wire \phy_ddio_dqdout[40] ;
wire \phy_ddio_dqdout[41] ;
wire \phy_ddio_dqdout[42] ;
wire \phy_ddio_dqdout[43] ;
wire \phy_ddio_dqdout[44] ;
wire \phy_ddio_dqdout[45] ;
wire \phy_ddio_dqdout[46] ;
wire \phy_ddio_dqdout[47] ;
wire \phy_ddio_dqdout[48] ;
wire \phy_ddio_dqdout[49] ;
wire \phy_ddio_dqdout[50] ;
wire \phy_ddio_dqdout[51] ;
wire \phy_ddio_dqdout[52] ;
wire \phy_ddio_dqdout[53] ;
wire \phy_ddio_dqdout[54] ;
wire \phy_ddio_dqdout[55] ;
wire \phy_ddio_dqdout[56] ;
wire \phy_ddio_dqdout[57] ;
wire \phy_ddio_dqdout[58] ;
wire \phy_ddio_dqdout[59] ;
wire \phy_ddio_dqdout[60] ;
wire \phy_ddio_dqdout[61] ;
wire \phy_ddio_dqdout[62] ;
wire \phy_ddio_dqdout[63] ;
wire \phy_ddio_dqdout[64] ;
wire \phy_ddio_dqdout[65] ;
wire \phy_ddio_dqdout[66] ;
wire \phy_ddio_dqdout[67] ;
wire \phy_ddio_dqdout[72] ;
wire \phy_ddio_dqdout[73] ;
wire \phy_ddio_dqdout[74] ;
wire \phy_ddio_dqdout[75] ;
wire \phy_ddio_dqdout[76] ;
wire \phy_ddio_dqdout[77] ;
wire \phy_ddio_dqdout[78] ;
wire \phy_ddio_dqdout[79] ;
wire \phy_ddio_dqdout[80] ;
wire \phy_ddio_dqdout[81] ;
wire \phy_ddio_dqdout[82] ;
wire \phy_ddio_dqdout[83] ;
wire \phy_ddio_dqdout[84] ;
wire \phy_ddio_dqdout[85] ;
wire \phy_ddio_dqdout[86] ;
wire \phy_ddio_dqdout[87] ;
wire \phy_ddio_dqdout[88] ;
wire \phy_ddio_dqdout[89] ;
wire \phy_ddio_dqdout[90] ;
wire \phy_ddio_dqdout[91] ;
wire \phy_ddio_dqdout[92] ;
wire \phy_ddio_dqdout[93] ;
wire \phy_ddio_dqdout[94] ;
wire \phy_ddio_dqdout[95] ;
wire \phy_ddio_dqdout[96] ;
wire \phy_ddio_dqdout[97] ;
wire \phy_ddio_dqdout[98] ;
wire \phy_ddio_dqdout[99] ;
wire \phy_ddio_dqdout[100] ;
wire \phy_ddio_dqdout[101] ;
wire \phy_ddio_dqdout[102] ;
wire \phy_ddio_dqdout[103] ;
wire \phy_ddio_dqdout[108] ;
wire \phy_ddio_dqdout[109] ;
wire \phy_ddio_dqdout[110] ;
wire \phy_ddio_dqdout[111] ;
wire \phy_ddio_dqdout[112] ;
wire \phy_ddio_dqdout[113] ;
wire \phy_ddio_dqdout[114] ;
wire \phy_ddio_dqdout[115] ;
wire \phy_ddio_dqdout[116] ;
wire \phy_ddio_dqdout[117] ;
wire \phy_ddio_dqdout[118] ;
wire \phy_ddio_dqdout[119] ;
wire \phy_ddio_dqdout[120] ;
wire \phy_ddio_dqdout[121] ;
wire \phy_ddio_dqdout[122] ;
wire \phy_ddio_dqdout[123] ;
wire \phy_ddio_dqdout[124] ;
wire \phy_ddio_dqdout[125] ;
wire \phy_ddio_dqdout[126] ;
wire \phy_ddio_dqdout[127] ;
wire \phy_ddio_dqdout[128] ;
wire \phy_ddio_dqdout[129] ;
wire \phy_ddio_dqdout[130] ;
wire \phy_ddio_dqdout[131] ;
wire \phy_ddio_dqdout[132] ;
wire \phy_ddio_dqdout[133] ;
wire \phy_ddio_dqdout[134] ;
wire \phy_ddio_dqdout[135] ;
wire \phy_ddio_dqdout[136] ;
wire \phy_ddio_dqdout[137] ;
wire \phy_ddio_dqdout[138] ;
wire \phy_ddio_dqdout[139] ;
wire \phy_ddio_dqoe[0] ;
wire \phy_ddio_dqoe[1] ;
wire \phy_ddio_dqoe[2] ;
wire \phy_ddio_dqoe[3] ;
wire \phy_ddio_dqoe[4] ;
wire \phy_ddio_dqoe[5] ;
wire \phy_ddio_dqoe[6] ;
wire \phy_ddio_dqoe[7] ;
wire \phy_ddio_dqoe[8] ;
wire \phy_ddio_dqoe[9] ;
wire \phy_ddio_dqoe[10] ;
wire \phy_ddio_dqoe[11] ;
wire \phy_ddio_dqoe[12] ;
wire \phy_ddio_dqoe[13] ;
wire \phy_ddio_dqoe[14] ;
wire \phy_ddio_dqoe[15] ;
wire \phy_ddio_dqoe[18] ;
wire \phy_ddio_dqoe[19] ;
wire \phy_ddio_dqoe[20] ;
wire \phy_ddio_dqoe[21] ;
wire \phy_ddio_dqoe[22] ;
wire \phy_ddio_dqoe[23] ;
wire \phy_ddio_dqoe[24] ;
wire \phy_ddio_dqoe[25] ;
wire \phy_ddio_dqoe[26] ;
wire \phy_ddio_dqoe[27] ;
wire \phy_ddio_dqoe[28] ;
wire \phy_ddio_dqoe[29] ;
wire \phy_ddio_dqoe[30] ;
wire \phy_ddio_dqoe[31] ;
wire \phy_ddio_dqoe[32] ;
wire \phy_ddio_dqoe[33] ;
wire \phy_ddio_dqoe[36] ;
wire \phy_ddio_dqoe[37] ;
wire \phy_ddio_dqoe[38] ;
wire \phy_ddio_dqoe[39] ;
wire \phy_ddio_dqoe[40] ;
wire \phy_ddio_dqoe[41] ;
wire \phy_ddio_dqoe[42] ;
wire \phy_ddio_dqoe[43] ;
wire \phy_ddio_dqoe[44] ;
wire \phy_ddio_dqoe[45] ;
wire \phy_ddio_dqoe[46] ;
wire \phy_ddio_dqoe[47] ;
wire \phy_ddio_dqoe[48] ;
wire \phy_ddio_dqoe[49] ;
wire \phy_ddio_dqoe[50] ;
wire \phy_ddio_dqoe[51] ;
wire \phy_ddio_dqoe[54] ;
wire \phy_ddio_dqoe[55] ;
wire \phy_ddio_dqoe[56] ;
wire \phy_ddio_dqoe[57] ;
wire \phy_ddio_dqoe[58] ;
wire \phy_ddio_dqoe[59] ;
wire \phy_ddio_dqoe[60] ;
wire \phy_ddio_dqoe[61] ;
wire \phy_ddio_dqoe[62] ;
wire \phy_ddio_dqoe[63] ;
wire \phy_ddio_dqoe[64] ;
wire \phy_ddio_dqoe[65] ;
wire \phy_ddio_dqoe[66] ;
wire \phy_ddio_dqoe[67] ;
wire \phy_ddio_dqoe[68] ;
wire \phy_ddio_dqoe[69] ;
wire \phy_ddio_dqs_dout[0] ;
wire \phy_ddio_dqs_dout[1] ;
wire \phy_ddio_dqs_dout[2] ;
wire \phy_ddio_dqs_dout[3] ;
wire \phy_ddio_dqs_dout[4] ;
wire \phy_ddio_dqs_dout[5] ;
wire \phy_ddio_dqs_dout[6] ;
wire \phy_ddio_dqs_dout[7] ;
wire \phy_ddio_dqs_dout[8] ;
wire \phy_ddio_dqs_dout[9] ;
wire \phy_ddio_dqs_dout[10] ;
wire \phy_ddio_dqs_dout[11] ;
wire \phy_ddio_dqs_dout[12] ;
wire \phy_ddio_dqs_dout[13] ;
wire \phy_ddio_dqs_dout[14] ;
wire \phy_ddio_dqs_dout[15] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[0] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[1] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[2] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[3] ;
wire \phy_ddio_dqslogic_aclr_pstamble[0] ;
wire \phy_ddio_dqslogic_aclr_pstamble[1] ;
wire \phy_ddio_dqslogic_aclr_pstamble[2] ;
wire \phy_ddio_dqslogic_aclr_pstamble[3] ;
wire \phy_ddio_dqslogic_dqsena[0] ;
wire \phy_ddio_dqslogic_dqsena[1] ;
wire \phy_ddio_dqslogic_dqsena[2] ;
wire \phy_ddio_dqslogic_dqsena[3] ;
wire \phy_ddio_dqslogic_dqsena[4] ;
wire \phy_ddio_dqslogic_dqsena[5] ;
wire \phy_ddio_dqslogic_dqsena[6] ;
wire \phy_ddio_dqslogic_dqsena[7] ;
wire \phy_ddio_dqslogic_fiforeset[0] ;
wire \phy_ddio_dqslogic_fiforeset[1] ;
wire \phy_ddio_dqslogic_fiforeset[2] ;
wire \phy_ddio_dqslogic_fiforeset[3] ;
wire \phy_ddio_dqslogic_incrdataen[0] ;
wire \phy_ddio_dqslogic_incrdataen[1] ;
wire \phy_ddio_dqslogic_incrdataen[2] ;
wire \phy_ddio_dqslogic_incrdataen[3] ;
wire \phy_ddio_dqslogic_incrdataen[4] ;
wire \phy_ddio_dqslogic_incrdataen[5] ;
wire \phy_ddio_dqslogic_incrdataen[6] ;
wire \phy_ddio_dqslogic_incrdataen[7] ;
wire \phy_ddio_dqslogic_incwrptr[0] ;
wire \phy_ddio_dqslogic_incwrptr[1] ;
wire \phy_ddio_dqslogic_incwrptr[2] ;
wire \phy_ddio_dqslogic_incwrptr[3] ;
wire \phy_ddio_dqslogic_incwrptr[4] ;
wire \phy_ddio_dqslogic_incwrptr[5] ;
wire \phy_ddio_dqslogic_incwrptr[6] ;
wire \phy_ddio_dqslogic_incwrptr[7] ;
wire \phy_ddio_dqslogic_oct[0] ;
wire \phy_ddio_dqslogic_oct[1] ;
wire \phy_ddio_dqslogic_oct[2] ;
wire \phy_ddio_dqslogic_oct[3] ;
wire \phy_ddio_dqslogic_oct[4] ;
wire \phy_ddio_dqslogic_oct[5] ;
wire \phy_ddio_dqslogic_oct[6] ;
wire \phy_ddio_dqslogic_oct[7] ;
wire \phy_ddio_dqslogic_readlatency[0] ;
wire \phy_ddio_dqslogic_readlatency[1] ;
wire \phy_ddio_dqslogic_readlatency[2] ;
wire \phy_ddio_dqslogic_readlatency[3] ;
wire \phy_ddio_dqslogic_readlatency[4] ;
wire \phy_ddio_dqslogic_readlatency[5] ;
wire \phy_ddio_dqslogic_readlatency[6] ;
wire \phy_ddio_dqslogic_readlatency[7] ;
wire \phy_ddio_dqslogic_readlatency[8] ;
wire \phy_ddio_dqslogic_readlatency[9] ;
wire \phy_ddio_dqslogic_readlatency[10] ;
wire \phy_ddio_dqslogic_readlatency[11] ;
wire \phy_ddio_dqslogic_readlatency[12] ;
wire \phy_ddio_dqslogic_readlatency[13] ;
wire \phy_ddio_dqslogic_readlatency[14] ;
wire \phy_ddio_dqslogic_readlatency[15] ;
wire \phy_ddio_dqslogic_readlatency[16] ;
wire \phy_ddio_dqslogic_readlatency[17] ;
wire \phy_ddio_dqslogic_readlatency[18] ;
wire \phy_ddio_dqslogic_readlatency[19] ;
wire \phy_ddio_dqs_oe[0] ;
wire \phy_ddio_dqs_oe[1] ;
wire \phy_ddio_dqs_oe[2] ;
wire \phy_ddio_dqs_oe[3] ;
wire \phy_ddio_dqs_oe[4] ;
wire \phy_ddio_dqs_oe[5] ;
wire \phy_ddio_dqs_oe[6] ;
wire \phy_ddio_dqs_oe[7] ;
wire \phy_ddio_odt[0] ;
wire \phy_ddio_odt[1] ;
wire \phy_ddio_odt[2] ;
wire \phy_ddio_odt[3] ;
wire \phy_ddio_ras_n[0] ;
wire \phy_ddio_ras_n[1] ;
wire \phy_ddio_ras_n[2] ;
wire \phy_ddio_ras_n[3] ;
wire \phy_ddio_reset_n[0] ;
wire \phy_ddio_reset_n[1] ;
wire \phy_ddio_reset_n[2] ;
wire \phy_ddio_reset_n[3] ;
wire \phy_ddio_we_n[0] ;
wire \phy_ddio_we_n[1] ;
wire \phy_ddio_we_n[2] ;
wire \phy_ddio_we_n[3] ;

wire [79:0] hphy_inst_AFIRDATA_bus;
wire [3:0] hphy_inst_AFIWLAT_bus;
wire [63:0] hphy_inst_PHYDDIOADDRDOUT_bus;
wire [11:0] hphy_inst_PHYDDIOBADOUT_bus;
wire [3:0] hphy_inst_PHYDDIOCASNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIOCKDOUT_bus;
wire [7:0] hphy_inst_PHYDDIOCKEDOUT_bus;
wire [7:0] hphy_inst_PHYDDIOCSNDOUT_bus;
wire [19:0] hphy_inst_PHYDDIODMDOUT_bus;
wire [179:0] hphy_inst_PHYDDIODQDOUT_bus;
wire [89:0] hphy_inst_PHYDDIODQOE_bus;
wire [19:0] hphy_inst_PHYDDIODQSDOUT_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICDQSENA_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICFIFORESET_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICOCT_bus;
wire [24:0] hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus;
wire [9:0] hphy_inst_PHYDDIODQSOE_bus;
wire [7:0] hphy_inst_PHYDDIOODTDOUT_bus;
wire [3:0] hphy_inst_PHYDDIORASNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIORESETNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIOWENDOUT_bus;

assign afi_rdata[0] = hphy_inst_AFIRDATA_bus[0];
assign afi_rdata[1] = hphy_inst_AFIRDATA_bus[1];
assign afi_rdata[2] = hphy_inst_AFIRDATA_bus[2];
assign afi_rdata[3] = hphy_inst_AFIRDATA_bus[3];
assign afi_rdata[4] = hphy_inst_AFIRDATA_bus[4];
assign afi_rdata[5] = hphy_inst_AFIRDATA_bus[5];
assign afi_rdata[6] = hphy_inst_AFIRDATA_bus[6];
assign afi_rdata[7] = hphy_inst_AFIRDATA_bus[7];
assign afi_rdata[8] = hphy_inst_AFIRDATA_bus[8];
assign afi_rdata[9] = hphy_inst_AFIRDATA_bus[9];
assign afi_rdata[10] = hphy_inst_AFIRDATA_bus[10];
assign afi_rdata[11] = hphy_inst_AFIRDATA_bus[11];
assign afi_rdata[12] = hphy_inst_AFIRDATA_bus[12];
assign afi_rdata[13] = hphy_inst_AFIRDATA_bus[13];
assign afi_rdata[14] = hphy_inst_AFIRDATA_bus[14];
assign afi_rdata[15] = hphy_inst_AFIRDATA_bus[15];
assign afi_rdata[16] = hphy_inst_AFIRDATA_bus[16];
assign afi_rdata[17] = hphy_inst_AFIRDATA_bus[17];
assign afi_rdata[18] = hphy_inst_AFIRDATA_bus[18];
assign afi_rdata[19] = hphy_inst_AFIRDATA_bus[19];
assign afi_rdata[20] = hphy_inst_AFIRDATA_bus[20];
assign afi_rdata[21] = hphy_inst_AFIRDATA_bus[21];
assign afi_rdata[22] = hphy_inst_AFIRDATA_bus[22];
assign afi_rdata[23] = hphy_inst_AFIRDATA_bus[23];
assign afi_rdata[24] = hphy_inst_AFIRDATA_bus[24];
assign afi_rdata[25] = hphy_inst_AFIRDATA_bus[25];
assign afi_rdata[26] = hphy_inst_AFIRDATA_bus[26];
assign afi_rdata[27] = hphy_inst_AFIRDATA_bus[27];
assign afi_rdata[28] = hphy_inst_AFIRDATA_bus[28];
assign afi_rdata[29] = hphy_inst_AFIRDATA_bus[29];
assign afi_rdata[30] = hphy_inst_AFIRDATA_bus[30];
assign afi_rdata[31] = hphy_inst_AFIRDATA_bus[31];
assign afi_rdata[32] = hphy_inst_AFIRDATA_bus[32];
assign afi_rdata[33] = hphy_inst_AFIRDATA_bus[33];
assign afi_rdata[34] = hphy_inst_AFIRDATA_bus[34];
assign afi_rdata[35] = hphy_inst_AFIRDATA_bus[35];
assign afi_rdata[36] = hphy_inst_AFIRDATA_bus[36];
assign afi_rdata[37] = hphy_inst_AFIRDATA_bus[37];
assign afi_rdata[38] = hphy_inst_AFIRDATA_bus[38];
assign afi_rdata[39] = hphy_inst_AFIRDATA_bus[39];
assign afi_rdata[40] = hphy_inst_AFIRDATA_bus[40];
assign afi_rdata[41] = hphy_inst_AFIRDATA_bus[41];
assign afi_rdata[42] = hphy_inst_AFIRDATA_bus[42];
assign afi_rdata[43] = hphy_inst_AFIRDATA_bus[43];
assign afi_rdata[44] = hphy_inst_AFIRDATA_bus[44];
assign afi_rdata[45] = hphy_inst_AFIRDATA_bus[45];
assign afi_rdata[46] = hphy_inst_AFIRDATA_bus[46];
assign afi_rdata[47] = hphy_inst_AFIRDATA_bus[47];
assign afi_rdata[48] = hphy_inst_AFIRDATA_bus[48];
assign afi_rdata[49] = hphy_inst_AFIRDATA_bus[49];
assign afi_rdata[50] = hphy_inst_AFIRDATA_bus[50];
assign afi_rdata[51] = hphy_inst_AFIRDATA_bus[51];
assign afi_rdata[52] = hphy_inst_AFIRDATA_bus[52];
assign afi_rdata[53] = hphy_inst_AFIRDATA_bus[53];
assign afi_rdata[54] = hphy_inst_AFIRDATA_bus[54];
assign afi_rdata[55] = hphy_inst_AFIRDATA_bus[55];
assign afi_rdata[56] = hphy_inst_AFIRDATA_bus[56];
assign afi_rdata[57] = hphy_inst_AFIRDATA_bus[57];
assign afi_rdata[58] = hphy_inst_AFIRDATA_bus[58];
assign afi_rdata[59] = hphy_inst_AFIRDATA_bus[59];
assign afi_rdata[60] = hphy_inst_AFIRDATA_bus[60];
assign afi_rdata[61] = hphy_inst_AFIRDATA_bus[61];
assign afi_rdata[62] = hphy_inst_AFIRDATA_bus[62];
assign afi_rdata[63] = hphy_inst_AFIRDATA_bus[63];
assign afi_rdata[64] = hphy_inst_AFIRDATA_bus[64];
assign afi_rdata[65] = hphy_inst_AFIRDATA_bus[65];
assign afi_rdata[66] = hphy_inst_AFIRDATA_bus[66];
assign afi_rdata[67] = hphy_inst_AFIRDATA_bus[67];
assign afi_rdata[68] = hphy_inst_AFIRDATA_bus[68];
assign afi_rdata[69] = hphy_inst_AFIRDATA_bus[69];
assign afi_rdata[70] = hphy_inst_AFIRDATA_bus[70];
assign afi_rdata[71] = hphy_inst_AFIRDATA_bus[71];
assign afi_rdata[72] = hphy_inst_AFIRDATA_bus[72];
assign afi_rdata[73] = hphy_inst_AFIRDATA_bus[73];
assign afi_rdata[74] = hphy_inst_AFIRDATA_bus[74];
assign afi_rdata[75] = hphy_inst_AFIRDATA_bus[75];
assign afi_rdata[76] = hphy_inst_AFIRDATA_bus[76];
assign afi_rdata[77] = hphy_inst_AFIRDATA_bus[77];
assign afi_rdata[78] = hphy_inst_AFIRDATA_bus[78];
assign afi_rdata[79] = hphy_inst_AFIRDATA_bus[79];

assign afi_wlat[0] = hphy_inst_AFIWLAT_bus[0];
assign afi_wlat[1] = hphy_inst_AFIWLAT_bus[1];
assign afi_wlat[2] = hphy_inst_AFIWLAT_bus[2];
assign afi_wlat[3] = hphy_inst_AFIWLAT_bus[3];

assign \phy_ddio_address[0]  = hphy_inst_PHYDDIOADDRDOUT_bus[0];
assign \phy_ddio_address[1]  = hphy_inst_PHYDDIOADDRDOUT_bus[1];
assign \phy_ddio_address[2]  = hphy_inst_PHYDDIOADDRDOUT_bus[2];
assign \phy_ddio_address[3]  = hphy_inst_PHYDDIOADDRDOUT_bus[3];
assign \phy_ddio_address[4]  = hphy_inst_PHYDDIOADDRDOUT_bus[4];
assign \phy_ddio_address[5]  = hphy_inst_PHYDDIOADDRDOUT_bus[5];
assign \phy_ddio_address[6]  = hphy_inst_PHYDDIOADDRDOUT_bus[6];
assign \phy_ddio_address[7]  = hphy_inst_PHYDDIOADDRDOUT_bus[7];
assign \phy_ddio_address[8]  = hphy_inst_PHYDDIOADDRDOUT_bus[8];
assign \phy_ddio_address[9]  = hphy_inst_PHYDDIOADDRDOUT_bus[9];
assign \phy_ddio_address[10]  = hphy_inst_PHYDDIOADDRDOUT_bus[10];
assign \phy_ddio_address[11]  = hphy_inst_PHYDDIOADDRDOUT_bus[11];
assign \phy_ddio_address[12]  = hphy_inst_PHYDDIOADDRDOUT_bus[12];
assign \phy_ddio_address[13]  = hphy_inst_PHYDDIOADDRDOUT_bus[13];
assign \phy_ddio_address[14]  = hphy_inst_PHYDDIOADDRDOUT_bus[14];
assign \phy_ddio_address[15]  = hphy_inst_PHYDDIOADDRDOUT_bus[15];
assign \phy_ddio_address[16]  = hphy_inst_PHYDDIOADDRDOUT_bus[16];
assign \phy_ddio_address[17]  = hphy_inst_PHYDDIOADDRDOUT_bus[17];
assign \phy_ddio_address[18]  = hphy_inst_PHYDDIOADDRDOUT_bus[18];
assign \phy_ddio_address[19]  = hphy_inst_PHYDDIOADDRDOUT_bus[19];
assign \phy_ddio_address[20]  = hphy_inst_PHYDDIOADDRDOUT_bus[20];
assign \phy_ddio_address[21]  = hphy_inst_PHYDDIOADDRDOUT_bus[21];
assign \phy_ddio_address[22]  = hphy_inst_PHYDDIOADDRDOUT_bus[22];
assign \phy_ddio_address[23]  = hphy_inst_PHYDDIOADDRDOUT_bus[23];
assign \phy_ddio_address[24]  = hphy_inst_PHYDDIOADDRDOUT_bus[24];
assign \phy_ddio_address[25]  = hphy_inst_PHYDDIOADDRDOUT_bus[25];
assign \phy_ddio_address[26]  = hphy_inst_PHYDDIOADDRDOUT_bus[26];
assign \phy_ddio_address[27]  = hphy_inst_PHYDDIOADDRDOUT_bus[27];
assign \phy_ddio_address[28]  = hphy_inst_PHYDDIOADDRDOUT_bus[28];
assign \phy_ddio_address[29]  = hphy_inst_PHYDDIOADDRDOUT_bus[29];
assign \phy_ddio_address[30]  = hphy_inst_PHYDDIOADDRDOUT_bus[30];
assign \phy_ddio_address[31]  = hphy_inst_PHYDDIOADDRDOUT_bus[31];
assign \phy_ddio_address[32]  = hphy_inst_PHYDDIOADDRDOUT_bus[32];
assign \phy_ddio_address[33]  = hphy_inst_PHYDDIOADDRDOUT_bus[33];
assign \phy_ddio_address[34]  = hphy_inst_PHYDDIOADDRDOUT_bus[34];
assign \phy_ddio_address[35]  = hphy_inst_PHYDDIOADDRDOUT_bus[35];
assign \phy_ddio_address[36]  = hphy_inst_PHYDDIOADDRDOUT_bus[36];
assign \phy_ddio_address[37]  = hphy_inst_PHYDDIOADDRDOUT_bus[37];
assign \phy_ddio_address[38]  = hphy_inst_PHYDDIOADDRDOUT_bus[38];
assign \phy_ddio_address[39]  = hphy_inst_PHYDDIOADDRDOUT_bus[39];
assign \phy_ddio_address[40]  = hphy_inst_PHYDDIOADDRDOUT_bus[40];
assign \phy_ddio_address[41]  = hphy_inst_PHYDDIOADDRDOUT_bus[41];
assign \phy_ddio_address[42]  = hphy_inst_PHYDDIOADDRDOUT_bus[42];
assign \phy_ddio_address[43]  = hphy_inst_PHYDDIOADDRDOUT_bus[43];
assign \phy_ddio_address[44]  = hphy_inst_PHYDDIOADDRDOUT_bus[44];
assign \phy_ddio_address[45]  = hphy_inst_PHYDDIOADDRDOUT_bus[45];
assign \phy_ddio_address[46]  = hphy_inst_PHYDDIOADDRDOUT_bus[46];
assign \phy_ddio_address[47]  = hphy_inst_PHYDDIOADDRDOUT_bus[47];
assign \phy_ddio_address[48]  = hphy_inst_PHYDDIOADDRDOUT_bus[48];
assign \phy_ddio_address[49]  = hphy_inst_PHYDDIOADDRDOUT_bus[49];
assign \phy_ddio_address[50]  = hphy_inst_PHYDDIOADDRDOUT_bus[50];
assign \phy_ddio_address[51]  = hphy_inst_PHYDDIOADDRDOUT_bus[51];
assign \phy_ddio_address[52]  = hphy_inst_PHYDDIOADDRDOUT_bus[52];
assign \phy_ddio_address[53]  = hphy_inst_PHYDDIOADDRDOUT_bus[53];
assign \phy_ddio_address[54]  = hphy_inst_PHYDDIOADDRDOUT_bus[54];
assign \phy_ddio_address[55]  = hphy_inst_PHYDDIOADDRDOUT_bus[55];
assign \phy_ddio_address[56]  = hphy_inst_PHYDDIOADDRDOUT_bus[56];
assign \phy_ddio_address[57]  = hphy_inst_PHYDDIOADDRDOUT_bus[57];
assign \phy_ddio_address[58]  = hphy_inst_PHYDDIOADDRDOUT_bus[58];
assign \phy_ddio_address[59]  = hphy_inst_PHYDDIOADDRDOUT_bus[59];

assign \phy_ddio_bank[0]  = hphy_inst_PHYDDIOBADOUT_bus[0];
assign \phy_ddio_bank[1]  = hphy_inst_PHYDDIOBADOUT_bus[1];
assign \phy_ddio_bank[2]  = hphy_inst_PHYDDIOBADOUT_bus[2];
assign \phy_ddio_bank[3]  = hphy_inst_PHYDDIOBADOUT_bus[3];
assign \phy_ddio_bank[4]  = hphy_inst_PHYDDIOBADOUT_bus[4];
assign \phy_ddio_bank[5]  = hphy_inst_PHYDDIOBADOUT_bus[5];
assign \phy_ddio_bank[6]  = hphy_inst_PHYDDIOBADOUT_bus[6];
assign \phy_ddio_bank[7]  = hphy_inst_PHYDDIOBADOUT_bus[7];
assign \phy_ddio_bank[8]  = hphy_inst_PHYDDIOBADOUT_bus[8];
assign \phy_ddio_bank[9]  = hphy_inst_PHYDDIOBADOUT_bus[9];
assign \phy_ddio_bank[10]  = hphy_inst_PHYDDIOBADOUT_bus[10];
assign \phy_ddio_bank[11]  = hphy_inst_PHYDDIOBADOUT_bus[11];

assign \phy_ddio_cas_n[0]  = hphy_inst_PHYDDIOCASNDOUT_bus[0];
assign \phy_ddio_cas_n[1]  = hphy_inst_PHYDDIOCASNDOUT_bus[1];
assign \phy_ddio_cas_n[2]  = hphy_inst_PHYDDIOCASNDOUT_bus[2];
assign \phy_ddio_cas_n[3]  = hphy_inst_PHYDDIOCASNDOUT_bus[3];

assign \phy_ddio_ck[0]  = hphy_inst_PHYDDIOCKDOUT_bus[0];
assign \phy_ddio_ck[1]  = hphy_inst_PHYDDIOCKDOUT_bus[1];

assign \phy_ddio_cke[0]  = hphy_inst_PHYDDIOCKEDOUT_bus[0];
assign \phy_ddio_cke[1]  = hphy_inst_PHYDDIOCKEDOUT_bus[1];
assign \phy_ddio_cke[2]  = hphy_inst_PHYDDIOCKEDOUT_bus[2];
assign \phy_ddio_cke[3]  = hphy_inst_PHYDDIOCKEDOUT_bus[3];

assign \phy_ddio_cs_n[0]  = hphy_inst_PHYDDIOCSNDOUT_bus[0];
assign \phy_ddio_cs_n[1]  = hphy_inst_PHYDDIOCSNDOUT_bus[1];
assign \phy_ddio_cs_n[2]  = hphy_inst_PHYDDIOCSNDOUT_bus[2];
assign \phy_ddio_cs_n[3]  = hphy_inst_PHYDDIOCSNDOUT_bus[3];

assign \phy_ddio_dmdout[0]  = hphy_inst_PHYDDIODMDOUT_bus[0];
assign \phy_ddio_dmdout[1]  = hphy_inst_PHYDDIODMDOUT_bus[1];
assign \phy_ddio_dmdout[2]  = hphy_inst_PHYDDIODMDOUT_bus[2];
assign \phy_ddio_dmdout[3]  = hphy_inst_PHYDDIODMDOUT_bus[3];
assign \phy_ddio_dmdout[4]  = hphy_inst_PHYDDIODMDOUT_bus[4];
assign \phy_ddio_dmdout[5]  = hphy_inst_PHYDDIODMDOUT_bus[5];
assign \phy_ddio_dmdout[6]  = hphy_inst_PHYDDIODMDOUT_bus[6];
assign \phy_ddio_dmdout[7]  = hphy_inst_PHYDDIODMDOUT_bus[7];
assign \phy_ddio_dmdout[8]  = hphy_inst_PHYDDIODMDOUT_bus[8];
assign \phy_ddio_dmdout[9]  = hphy_inst_PHYDDIODMDOUT_bus[9];
assign \phy_ddio_dmdout[10]  = hphy_inst_PHYDDIODMDOUT_bus[10];
assign \phy_ddio_dmdout[11]  = hphy_inst_PHYDDIODMDOUT_bus[11];
assign \phy_ddio_dmdout[12]  = hphy_inst_PHYDDIODMDOUT_bus[12];
assign \phy_ddio_dmdout[13]  = hphy_inst_PHYDDIODMDOUT_bus[13];
assign \phy_ddio_dmdout[14]  = hphy_inst_PHYDDIODMDOUT_bus[14];
assign \phy_ddio_dmdout[15]  = hphy_inst_PHYDDIODMDOUT_bus[15];

assign \phy_ddio_dqdout[0]  = hphy_inst_PHYDDIODQDOUT_bus[0];
assign \phy_ddio_dqdout[1]  = hphy_inst_PHYDDIODQDOUT_bus[1];
assign \phy_ddio_dqdout[2]  = hphy_inst_PHYDDIODQDOUT_bus[2];
assign \phy_ddio_dqdout[3]  = hphy_inst_PHYDDIODQDOUT_bus[3];
assign \phy_ddio_dqdout[4]  = hphy_inst_PHYDDIODQDOUT_bus[4];
assign \phy_ddio_dqdout[5]  = hphy_inst_PHYDDIODQDOUT_bus[5];
assign \phy_ddio_dqdout[6]  = hphy_inst_PHYDDIODQDOUT_bus[6];
assign \phy_ddio_dqdout[7]  = hphy_inst_PHYDDIODQDOUT_bus[7];
assign \phy_ddio_dqdout[8]  = hphy_inst_PHYDDIODQDOUT_bus[8];
assign \phy_ddio_dqdout[9]  = hphy_inst_PHYDDIODQDOUT_bus[9];
assign \phy_ddio_dqdout[10]  = hphy_inst_PHYDDIODQDOUT_bus[10];
assign \phy_ddio_dqdout[11]  = hphy_inst_PHYDDIODQDOUT_bus[11];
assign \phy_ddio_dqdout[12]  = hphy_inst_PHYDDIODQDOUT_bus[12];
assign \phy_ddio_dqdout[13]  = hphy_inst_PHYDDIODQDOUT_bus[13];
assign \phy_ddio_dqdout[14]  = hphy_inst_PHYDDIODQDOUT_bus[14];
assign \phy_ddio_dqdout[15]  = hphy_inst_PHYDDIODQDOUT_bus[15];
assign \phy_ddio_dqdout[16]  = hphy_inst_PHYDDIODQDOUT_bus[16];
assign \phy_ddio_dqdout[17]  = hphy_inst_PHYDDIODQDOUT_bus[17];
assign \phy_ddio_dqdout[18]  = hphy_inst_PHYDDIODQDOUT_bus[18];
assign \phy_ddio_dqdout[19]  = hphy_inst_PHYDDIODQDOUT_bus[19];
assign \phy_ddio_dqdout[20]  = hphy_inst_PHYDDIODQDOUT_bus[20];
assign \phy_ddio_dqdout[21]  = hphy_inst_PHYDDIODQDOUT_bus[21];
assign \phy_ddio_dqdout[22]  = hphy_inst_PHYDDIODQDOUT_bus[22];
assign \phy_ddio_dqdout[23]  = hphy_inst_PHYDDIODQDOUT_bus[23];
assign \phy_ddio_dqdout[24]  = hphy_inst_PHYDDIODQDOUT_bus[24];
assign \phy_ddio_dqdout[25]  = hphy_inst_PHYDDIODQDOUT_bus[25];
assign \phy_ddio_dqdout[26]  = hphy_inst_PHYDDIODQDOUT_bus[26];
assign \phy_ddio_dqdout[27]  = hphy_inst_PHYDDIODQDOUT_bus[27];
assign \phy_ddio_dqdout[28]  = hphy_inst_PHYDDIODQDOUT_bus[28];
assign \phy_ddio_dqdout[29]  = hphy_inst_PHYDDIODQDOUT_bus[29];
assign \phy_ddio_dqdout[30]  = hphy_inst_PHYDDIODQDOUT_bus[30];
assign \phy_ddio_dqdout[31]  = hphy_inst_PHYDDIODQDOUT_bus[31];
assign \phy_ddio_dqdout[36]  = hphy_inst_PHYDDIODQDOUT_bus[36];
assign \phy_ddio_dqdout[37]  = hphy_inst_PHYDDIODQDOUT_bus[37];
assign \phy_ddio_dqdout[38]  = hphy_inst_PHYDDIODQDOUT_bus[38];
assign \phy_ddio_dqdout[39]  = hphy_inst_PHYDDIODQDOUT_bus[39];
assign \phy_ddio_dqdout[40]  = hphy_inst_PHYDDIODQDOUT_bus[40];
assign \phy_ddio_dqdout[41]  = hphy_inst_PHYDDIODQDOUT_bus[41];
assign \phy_ddio_dqdout[42]  = hphy_inst_PHYDDIODQDOUT_bus[42];
assign \phy_ddio_dqdout[43]  = hphy_inst_PHYDDIODQDOUT_bus[43];
assign \phy_ddio_dqdout[44]  = hphy_inst_PHYDDIODQDOUT_bus[44];
assign \phy_ddio_dqdout[45]  = hphy_inst_PHYDDIODQDOUT_bus[45];
assign \phy_ddio_dqdout[46]  = hphy_inst_PHYDDIODQDOUT_bus[46];
assign \phy_ddio_dqdout[47]  = hphy_inst_PHYDDIODQDOUT_bus[47];
assign \phy_ddio_dqdout[48]  = hphy_inst_PHYDDIODQDOUT_bus[48];
assign \phy_ddio_dqdout[49]  = hphy_inst_PHYDDIODQDOUT_bus[49];
assign \phy_ddio_dqdout[50]  = hphy_inst_PHYDDIODQDOUT_bus[50];
assign \phy_ddio_dqdout[51]  = hphy_inst_PHYDDIODQDOUT_bus[51];
assign \phy_ddio_dqdout[52]  = hphy_inst_PHYDDIODQDOUT_bus[52];
assign \phy_ddio_dqdout[53]  = hphy_inst_PHYDDIODQDOUT_bus[53];
assign \phy_ddio_dqdout[54]  = hphy_inst_PHYDDIODQDOUT_bus[54];
assign \phy_ddio_dqdout[55]  = hphy_inst_PHYDDIODQDOUT_bus[55];
assign \phy_ddio_dqdout[56]  = hphy_inst_PHYDDIODQDOUT_bus[56];
assign \phy_ddio_dqdout[57]  = hphy_inst_PHYDDIODQDOUT_bus[57];
assign \phy_ddio_dqdout[58]  = hphy_inst_PHYDDIODQDOUT_bus[58];
assign \phy_ddio_dqdout[59]  = hphy_inst_PHYDDIODQDOUT_bus[59];
assign \phy_ddio_dqdout[60]  = hphy_inst_PHYDDIODQDOUT_bus[60];
assign \phy_ddio_dqdout[61]  = hphy_inst_PHYDDIODQDOUT_bus[61];
assign \phy_ddio_dqdout[62]  = hphy_inst_PHYDDIODQDOUT_bus[62];
assign \phy_ddio_dqdout[63]  = hphy_inst_PHYDDIODQDOUT_bus[63];
assign \phy_ddio_dqdout[64]  = hphy_inst_PHYDDIODQDOUT_bus[64];
assign \phy_ddio_dqdout[65]  = hphy_inst_PHYDDIODQDOUT_bus[65];
assign \phy_ddio_dqdout[66]  = hphy_inst_PHYDDIODQDOUT_bus[66];
assign \phy_ddio_dqdout[67]  = hphy_inst_PHYDDIODQDOUT_bus[67];
assign \phy_ddio_dqdout[72]  = hphy_inst_PHYDDIODQDOUT_bus[72];
assign \phy_ddio_dqdout[73]  = hphy_inst_PHYDDIODQDOUT_bus[73];
assign \phy_ddio_dqdout[74]  = hphy_inst_PHYDDIODQDOUT_bus[74];
assign \phy_ddio_dqdout[75]  = hphy_inst_PHYDDIODQDOUT_bus[75];
assign \phy_ddio_dqdout[76]  = hphy_inst_PHYDDIODQDOUT_bus[76];
assign \phy_ddio_dqdout[77]  = hphy_inst_PHYDDIODQDOUT_bus[77];
assign \phy_ddio_dqdout[78]  = hphy_inst_PHYDDIODQDOUT_bus[78];
assign \phy_ddio_dqdout[79]  = hphy_inst_PHYDDIODQDOUT_bus[79];
assign \phy_ddio_dqdout[80]  = hphy_inst_PHYDDIODQDOUT_bus[80];
assign \phy_ddio_dqdout[81]  = hphy_inst_PHYDDIODQDOUT_bus[81];
assign \phy_ddio_dqdout[82]  = hphy_inst_PHYDDIODQDOUT_bus[82];
assign \phy_ddio_dqdout[83]  = hphy_inst_PHYDDIODQDOUT_bus[83];
assign \phy_ddio_dqdout[84]  = hphy_inst_PHYDDIODQDOUT_bus[84];
assign \phy_ddio_dqdout[85]  = hphy_inst_PHYDDIODQDOUT_bus[85];
assign \phy_ddio_dqdout[86]  = hphy_inst_PHYDDIODQDOUT_bus[86];
assign \phy_ddio_dqdout[87]  = hphy_inst_PHYDDIODQDOUT_bus[87];
assign \phy_ddio_dqdout[88]  = hphy_inst_PHYDDIODQDOUT_bus[88];
assign \phy_ddio_dqdout[89]  = hphy_inst_PHYDDIODQDOUT_bus[89];
assign \phy_ddio_dqdout[90]  = hphy_inst_PHYDDIODQDOUT_bus[90];
assign \phy_ddio_dqdout[91]  = hphy_inst_PHYDDIODQDOUT_bus[91];
assign \phy_ddio_dqdout[92]  = hphy_inst_PHYDDIODQDOUT_bus[92];
assign \phy_ddio_dqdout[93]  = hphy_inst_PHYDDIODQDOUT_bus[93];
assign \phy_ddio_dqdout[94]  = hphy_inst_PHYDDIODQDOUT_bus[94];
assign \phy_ddio_dqdout[95]  = hphy_inst_PHYDDIODQDOUT_bus[95];
assign \phy_ddio_dqdout[96]  = hphy_inst_PHYDDIODQDOUT_bus[96];
assign \phy_ddio_dqdout[97]  = hphy_inst_PHYDDIODQDOUT_bus[97];
assign \phy_ddio_dqdout[98]  = hphy_inst_PHYDDIODQDOUT_bus[98];
assign \phy_ddio_dqdout[99]  = hphy_inst_PHYDDIODQDOUT_bus[99];
assign \phy_ddio_dqdout[100]  = hphy_inst_PHYDDIODQDOUT_bus[100];
assign \phy_ddio_dqdout[101]  = hphy_inst_PHYDDIODQDOUT_bus[101];
assign \phy_ddio_dqdout[102]  = hphy_inst_PHYDDIODQDOUT_bus[102];
assign \phy_ddio_dqdout[103]  = hphy_inst_PHYDDIODQDOUT_bus[103];
assign \phy_ddio_dqdout[108]  = hphy_inst_PHYDDIODQDOUT_bus[108];
assign \phy_ddio_dqdout[109]  = hphy_inst_PHYDDIODQDOUT_bus[109];
assign \phy_ddio_dqdout[110]  = hphy_inst_PHYDDIODQDOUT_bus[110];
assign \phy_ddio_dqdout[111]  = hphy_inst_PHYDDIODQDOUT_bus[111];
assign \phy_ddio_dqdout[112]  = hphy_inst_PHYDDIODQDOUT_bus[112];
assign \phy_ddio_dqdout[113]  = hphy_inst_PHYDDIODQDOUT_bus[113];
assign \phy_ddio_dqdout[114]  = hphy_inst_PHYDDIODQDOUT_bus[114];
assign \phy_ddio_dqdout[115]  = hphy_inst_PHYDDIODQDOUT_bus[115];
assign \phy_ddio_dqdout[116]  = hphy_inst_PHYDDIODQDOUT_bus[116];
assign \phy_ddio_dqdout[117]  = hphy_inst_PHYDDIODQDOUT_bus[117];
assign \phy_ddio_dqdout[118]  = hphy_inst_PHYDDIODQDOUT_bus[118];
assign \phy_ddio_dqdout[119]  = hphy_inst_PHYDDIODQDOUT_bus[119];
assign \phy_ddio_dqdout[120]  = hphy_inst_PHYDDIODQDOUT_bus[120];
assign \phy_ddio_dqdout[121]  = hphy_inst_PHYDDIODQDOUT_bus[121];
assign \phy_ddio_dqdout[122]  = hphy_inst_PHYDDIODQDOUT_bus[122];
assign \phy_ddio_dqdout[123]  = hphy_inst_PHYDDIODQDOUT_bus[123];
assign \phy_ddio_dqdout[124]  = hphy_inst_PHYDDIODQDOUT_bus[124];
assign \phy_ddio_dqdout[125]  = hphy_inst_PHYDDIODQDOUT_bus[125];
assign \phy_ddio_dqdout[126]  = hphy_inst_PHYDDIODQDOUT_bus[126];
assign \phy_ddio_dqdout[127]  = hphy_inst_PHYDDIODQDOUT_bus[127];
assign \phy_ddio_dqdout[128]  = hphy_inst_PHYDDIODQDOUT_bus[128];
assign \phy_ddio_dqdout[129]  = hphy_inst_PHYDDIODQDOUT_bus[129];
assign \phy_ddio_dqdout[130]  = hphy_inst_PHYDDIODQDOUT_bus[130];
assign \phy_ddio_dqdout[131]  = hphy_inst_PHYDDIODQDOUT_bus[131];
assign \phy_ddio_dqdout[132]  = hphy_inst_PHYDDIODQDOUT_bus[132];
assign \phy_ddio_dqdout[133]  = hphy_inst_PHYDDIODQDOUT_bus[133];
assign \phy_ddio_dqdout[134]  = hphy_inst_PHYDDIODQDOUT_bus[134];
assign \phy_ddio_dqdout[135]  = hphy_inst_PHYDDIODQDOUT_bus[135];
assign \phy_ddio_dqdout[136]  = hphy_inst_PHYDDIODQDOUT_bus[136];
assign \phy_ddio_dqdout[137]  = hphy_inst_PHYDDIODQDOUT_bus[137];
assign \phy_ddio_dqdout[138]  = hphy_inst_PHYDDIODQDOUT_bus[138];
assign \phy_ddio_dqdout[139]  = hphy_inst_PHYDDIODQDOUT_bus[139];

assign \phy_ddio_dqoe[0]  = hphy_inst_PHYDDIODQOE_bus[0];
assign \phy_ddio_dqoe[1]  = hphy_inst_PHYDDIODQOE_bus[1];
assign \phy_ddio_dqoe[2]  = hphy_inst_PHYDDIODQOE_bus[2];
assign \phy_ddio_dqoe[3]  = hphy_inst_PHYDDIODQOE_bus[3];
assign \phy_ddio_dqoe[4]  = hphy_inst_PHYDDIODQOE_bus[4];
assign \phy_ddio_dqoe[5]  = hphy_inst_PHYDDIODQOE_bus[5];
assign \phy_ddio_dqoe[6]  = hphy_inst_PHYDDIODQOE_bus[6];
assign \phy_ddio_dqoe[7]  = hphy_inst_PHYDDIODQOE_bus[7];
assign \phy_ddio_dqoe[8]  = hphy_inst_PHYDDIODQOE_bus[8];
assign \phy_ddio_dqoe[9]  = hphy_inst_PHYDDIODQOE_bus[9];
assign \phy_ddio_dqoe[10]  = hphy_inst_PHYDDIODQOE_bus[10];
assign \phy_ddio_dqoe[11]  = hphy_inst_PHYDDIODQOE_bus[11];
assign \phy_ddio_dqoe[12]  = hphy_inst_PHYDDIODQOE_bus[12];
assign \phy_ddio_dqoe[13]  = hphy_inst_PHYDDIODQOE_bus[13];
assign \phy_ddio_dqoe[14]  = hphy_inst_PHYDDIODQOE_bus[14];
assign \phy_ddio_dqoe[15]  = hphy_inst_PHYDDIODQOE_bus[15];
assign \phy_ddio_dqoe[18]  = hphy_inst_PHYDDIODQOE_bus[18];
assign \phy_ddio_dqoe[19]  = hphy_inst_PHYDDIODQOE_bus[19];
assign \phy_ddio_dqoe[20]  = hphy_inst_PHYDDIODQOE_bus[20];
assign \phy_ddio_dqoe[21]  = hphy_inst_PHYDDIODQOE_bus[21];
assign \phy_ddio_dqoe[22]  = hphy_inst_PHYDDIODQOE_bus[22];
assign \phy_ddio_dqoe[23]  = hphy_inst_PHYDDIODQOE_bus[23];
assign \phy_ddio_dqoe[24]  = hphy_inst_PHYDDIODQOE_bus[24];
assign \phy_ddio_dqoe[25]  = hphy_inst_PHYDDIODQOE_bus[25];
assign \phy_ddio_dqoe[26]  = hphy_inst_PHYDDIODQOE_bus[26];
assign \phy_ddio_dqoe[27]  = hphy_inst_PHYDDIODQOE_bus[27];
assign \phy_ddio_dqoe[28]  = hphy_inst_PHYDDIODQOE_bus[28];
assign \phy_ddio_dqoe[29]  = hphy_inst_PHYDDIODQOE_bus[29];
assign \phy_ddio_dqoe[30]  = hphy_inst_PHYDDIODQOE_bus[30];
assign \phy_ddio_dqoe[31]  = hphy_inst_PHYDDIODQOE_bus[31];
assign \phy_ddio_dqoe[32]  = hphy_inst_PHYDDIODQOE_bus[32];
assign \phy_ddio_dqoe[33]  = hphy_inst_PHYDDIODQOE_bus[33];
assign \phy_ddio_dqoe[36]  = hphy_inst_PHYDDIODQOE_bus[36];
assign \phy_ddio_dqoe[37]  = hphy_inst_PHYDDIODQOE_bus[37];
assign \phy_ddio_dqoe[38]  = hphy_inst_PHYDDIODQOE_bus[38];
assign \phy_ddio_dqoe[39]  = hphy_inst_PHYDDIODQOE_bus[39];
assign \phy_ddio_dqoe[40]  = hphy_inst_PHYDDIODQOE_bus[40];
assign \phy_ddio_dqoe[41]  = hphy_inst_PHYDDIODQOE_bus[41];
assign \phy_ddio_dqoe[42]  = hphy_inst_PHYDDIODQOE_bus[42];
assign \phy_ddio_dqoe[43]  = hphy_inst_PHYDDIODQOE_bus[43];
assign \phy_ddio_dqoe[44]  = hphy_inst_PHYDDIODQOE_bus[44];
assign \phy_ddio_dqoe[45]  = hphy_inst_PHYDDIODQOE_bus[45];
assign \phy_ddio_dqoe[46]  = hphy_inst_PHYDDIODQOE_bus[46];
assign \phy_ddio_dqoe[47]  = hphy_inst_PHYDDIODQOE_bus[47];
assign \phy_ddio_dqoe[48]  = hphy_inst_PHYDDIODQOE_bus[48];
assign \phy_ddio_dqoe[49]  = hphy_inst_PHYDDIODQOE_bus[49];
assign \phy_ddio_dqoe[50]  = hphy_inst_PHYDDIODQOE_bus[50];
assign \phy_ddio_dqoe[51]  = hphy_inst_PHYDDIODQOE_bus[51];
assign \phy_ddio_dqoe[54]  = hphy_inst_PHYDDIODQOE_bus[54];
assign \phy_ddio_dqoe[55]  = hphy_inst_PHYDDIODQOE_bus[55];
assign \phy_ddio_dqoe[56]  = hphy_inst_PHYDDIODQOE_bus[56];
assign \phy_ddio_dqoe[57]  = hphy_inst_PHYDDIODQOE_bus[57];
assign \phy_ddio_dqoe[58]  = hphy_inst_PHYDDIODQOE_bus[58];
assign \phy_ddio_dqoe[59]  = hphy_inst_PHYDDIODQOE_bus[59];
assign \phy_ddio_dqoe[60]  = hphy_inst_PHYDDIODQOE_bus[60];
assign \phy_ddio_dqoe[61]  = hphy_inst_PHYDDIODQOE_bus[61];
assign \phy_ddio_dqoe[62]  = hphy_inst_PHYDDIODQOE_bus[62];
assign \phy_ddio_dqoe[63]  = hphy_inst_PHYDDIODQOE_bus[63];
assign \phy_ddio_dqoe[64]  = hphy_inst_PHYDDIODQOE_bus[64];
assign \phy_ddio_dqoe[65]  = hphy_inst_PHYDDIODQOE_bus[65];
assign \phy_ddio_dqoe[66]  = hphy_inst_PHYDDIODQOE_bus[66];
assign \phy_ddio_dqoe[67]  = hphy_inst_PHYDDIODQOE_bus[67];
assign \phy_ddio_dqoe[68]  = hphy_inst_PHYDDIODQOE_bus[68];
assign \phy_ddio_dqoe[69]  = hphy_inst_PHYDDIODQOE_bus[69];

assign \phy_ddio_dqs_dout[0]  = hphy_inst_PHYDDIODQSDOUT_bus[0];
assign \phy_ddio_dqs_dout[1]  = hphy_inst_PHYDDIODQSDOUT_bus[1];
assign \phy_ddio_dqs_dout[2]  = hphy_inst_PHYDDIODQSDOUT_bus[2];
assign \phy_ddio_dqs_dout[3]  = hphy_inst_PHYDDIODQSDOUT_bus[3];
assign \phy_ddio_dqs_dout[4]  = hphy_inst_PHYDDIODQSDOUT_bus[4];
assign \phy_ddio_dqs_dout[5]  = hphy_inst_PHYDDIODQSDOUT_bus[5];
assign \phy_ddio_dqs_dout[6]  = hphy_inst_PHYDDIODQSDOUT_bus[6];
assign \phy_ddio_dqs_dout[7]  = hphy_inst_PHYDDIODQSDOUT_bus[7];
assign \phy_ddio_dqs_dout[8]  = hphy_inst_PHYDDIODQSDOUT_bus[8];
assign \phy_ddio_dqs_dout[9]  = hphy_inst_PHYDDIODQSDOUT_bus[9];
assign \phy_ddio_dqs_dout[10]  = hphy_inst_PHYDDIODQSDOUT_bus[10];
assign \phy_ddio_dqs_dout[11]  = hphy_inst_PHYDDIODQSDOUT_bus[11];
assign \phy_ddio_dqs_dout[12]  = hphy_inst_PHYDDIODQSDOUT_bus[12];
assign \phy_ddio_dqs_dout[13]  = hphy_inst_PHYDDIODQSDOUT_bus[13];
assign \phy_ddio_dqs_dout[14]  = hphy_inst_PHYDDIODQSDOUT_bus[14];
assign \phy_ddio_dqs_dout[15]  = hphy_inst_PHYDDIODQSDOUT_bus[15];

assign \phy_ddio_dqslogic_aclr_fifoctrl[0]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[0];
assign \phy_ddio_dqslogic_aclr_fifoctrl[1]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[1];
assign \phy_ddio_dqslogic_aclr_fifoctrl[2]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[2];
assign \phy_ddio_dqslogic_aclr_fifoctrl[3]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[3];

assign \phy_ddio_dqslogic_aclr_pstamble[0]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[0];
assign \phy_ddio_dqslogic_aclr_pstamble[1]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[1];
assign \phy_ddio_dqslogic_aclr_pstamble[2]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[2];
assign \phy_ddio_dqslogic_aclr_pstamble[3]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[3];

assign \phy_ddio_dqslogic_dqsena[0]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[0];
assign \phy_ddio_dqslogic_dqsena[1]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[1];
assign \phy_ddio_dqslogic_dqsena[2]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[2];
assign \phy_ddio_dqslogic_dqsena[3]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[3];
assign \phy_ddio_dqslogic_dqsena[4]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[4];
assign \phy_ddio_dqslogic_dqsena[5]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[5];
assign \phy_ddio_dqslogic_dqsena[6]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[6];
assign \phy_ddio_dqslogic_dqsena[7]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[7];

assign \phy_ddio_dqslogic_fiforeset[0]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[0];
assign \phy_ddio_dqslogic_fiforeset[1]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[1];
assign \phy_ddio_dqslogic_fiforeset[2]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[2];
assign \phy_ddio_dqslogic_fiforeset[3]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[3];

assign \phy_ddio_dqslogic_incrdataen[0]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[0];
assign \phy_ddio_dqslogic_incrdataen[1]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[1];
assign \phy_ddio_dqslogic_incrdataen[2]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[2];
assign \phy_ddio_dqslogic_incrdataen[3]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[3];
assign \phy_ddio_dqslogic_incrdataen[4]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[4];
assign \phy_ddio_dqslogic_incrdataen[5]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[5];
assign \phy_ddio_dqslogic_incrdataen[6]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[6];
assign \phy_ddio_dqslogic_incrdataen[7]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[7];

assign \phy_ddio_dqslogic_incwrptr[0]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[0];
assign \phy_ddio_dqslogic_incwrptr[1]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[1];
assign \phy_ddio_dqslogic_incwrptr[2]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[2];
assign \phy_ddio_dqslogic_incwrptr[3]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[3];
assign \phy_ddio_dqslogic_incwrptr[4]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[4];
assign \phy_ddio_dqslogic_incwrptr[5]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[5];
assign \phy_ddio_dqslogic_incwrptr[6]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[6];
assign \phy_ddio_dqslogic_incwrptr[7]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[7];

assign \phy_ddio_dqslogic_oct[0]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[0];
assign \phy_ddio_dqslogic_oct[1]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[1];
assign \phy_ddio_dqslogic_oct[2]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[2];
assign \phy_ddio_dqslogic_oct[3]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[3];
assign \phy_ddio_dqslogic_oct[4]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[4];
assign \phy_ddio_dqslogic_oct[5]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[5];
assign \phy_ddio_dqslogic_oct[6]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[6];
assign \phy_ddio_dqslogic_oct[7]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[7];

assign \phy_ddio_dqslogic_readlatency[0]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[0];
assign \phy_ddio_dqslogic_readlatency[1]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[1];
assign \phy_ddio_dqslogic_readlatency[2]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[2];
assign \phy_ddio_dqslogic_readlatency[3]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[3];
assign \phy_ddio_dqslogic_readlatency[4]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[4];
assign \phy_ddio_dqslogic_readlatency[5]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[5];
assign \phy_ddio_dqslogic_readlatency[6]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[6];
assign \phy_ddio_dqslogic_readlatency[7]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[7];
assign \phy_ddio_dqslogic_readlatency[8]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[8];
assign \phy_ddio_dqslogic_readlatency[9]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[9];
assign \phy_ddio_dqslogic_readlatency[10]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[10];
assign \phy_ddio_dqslogic_readlatency[11]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[11];
assign \phy_ddio_dqslogic_readlatency[12]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[12];
assign \phy_ddio_dqslogic_readlatency[13]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[13];
assign \phy_ddio_dqslogic_readlatency[14]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[14];
assign \phy_ddio_dqslogic_readlatency[15]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[15];
assign \phy_ddio_dqslogic_readlatency[16]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[16];
assign \phy_ddio_dqslogic_readlatency[17]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[17];
assign \phy_ddio_dqslogic_readlatency[18]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[18];
assign \phy_ddio_dqslogic_readlatency[19]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[19];

assign \phy_ddio_dqs_oe[0]  = hphy_inst_PHYDDIODQSOE_bus[0];
assign \phy_ddio_dqs_oe[1]  = hphy_inst_PHYDDIODQSOE_bus[1];
assign \phy_ddio_dqs_oe[2]  = hphy_inst_PHYDDIODQSOE_bus[2];
assign \phy_ddio_dqs_oe[3]  = hphy_inst_PHYDDIODQSOE_bus[3];
assign \phy_ddio_dqs_oe[4]  = hphy_inst_PHYDDIODQSOE_bus[4];
assign \phy_ddio_dqs_oe[5]  = hphy_inst_PHYDDIODQSOE_bus[5];
assign \phy_ddio_dqs_oe[6]  = hphy_inst_PHYDDIODQSOE_bus[6];
assign \phy_ddio_dqs_oe[7]  = hphy_inst_PHYDDIODQSOE_bus[7];

assign \phy_ddio_odt[0]  = hphy_inst_PHYDDIOODTDOUT_bus[0];
assign \phy_ddio_odt[1]  = hphy_inst_PHYDDIOODTDOUT_bus[1];
assign \phy_ddio_odt[2]  = hphy_inst_PHYDDIOODTDOUT_bus[2];
assign \phy_ddio_odt[3]  = hphy_inst_PHYDDIOODTDOUT_bus[3];

assign \phy_ddio_ras_n[0]  = hphy_inst_PHYDDIORASNDOUT_bus[0];
assign \phy_ddio_ras_n[1]  = hphy_inst_PHYDDIORASNDOUT_bus[1];
assign \phy_ddio_ras_n[2]  = hphy_inst_PHYDDIORASNDOUT_bus[2];
assign \phy_ddio_ras_n[3]  = hphy_inst_PHYDDIORASNDOUT_bus[3];

assign \phy_ddio_reset_n[0]  = hphy_inst_PHYDDIORESETNDOUT_bus[0];
assign \phy_ddio_reset_n[1]  = hphy_inst_PHYDDIORESETNDOUT_bus[1];
assign \phy_ddio_reset_n[2]  = hphy_inst_PHYDDIORESETNDOUT_bus[2];
assign \phy_ddio_reset_n[3]  = hphy_inst_PHYDDIORESETNDOUT_bus[3];

assign \phy_ddio_we_n[0]  = hphy_inst_PHYDDIOWENDOUT_bus[0];
assign \phy_ddio_we_n[1]  = hphy_inst_PHYDDIOWENDOUT_bus[1];
assign \phy_ddio_we_n[2]  = hphy_inst_PHYDDIOWENDOUT_bus[2];
assign \phy_ddio_we_n[3]  = hphy_inst_PHYDDIOWENDOUT_bus[3];

Computer_System_hps_sdram_p0_acv_hard_io_pads uio_pads(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.phy_ddio_address_0(\phy_ddio_address[0] ),
	.phy_ddio_address_1(\phy_ddio_address[1] ),
	.phy_ddio_address_2(\phy_ddio_address[2] ),
	.phy_ddio_address_3(\phy_ddio_address[3] ),
	.phy_ddio_address_4(\phy_ddio_address[4] ),
	.phy_ddio_address_5(\phy_ddio_address[5] ),
	.phy_ddio_address_6(\phy_ddio_address[6] ),
	.phy_ddio_address_7(\phy_ddio_address[7] ),
	.phy_ddio_address_8(\phy_ddio_address[8] ),
	.phy_ddio_address_9(\phy_ddio_address[9] ),
	.phy_ddio_address_10(\phy_ddio_address[10] ),
	.phy_ddio_address_11(\phy_ddio_address[11] ),
	.phy_ddio_address_12(\phy_ddio_address[12] ),
	.phy_ddio_address_13(\phy_ddio_address[13] ),
	.phy_ddio_address_14(\phy_ddio_address[14] ),
	.phy_ddio_address_15(\phy_ddio_address[15] ),
	.phy_ddio_address_16(\phy_ddio_address[16] ),
	.phy_ddio_address_17(\phy_ddio_address[17] ),
	.phy_ddio_address_18(\phy_ddio_address[18] ),
	.phy_ddio_address_19(\phy_ddio_address[19] ),
	.phy_ddio_address_20(\phy_ddio_address[20] ),
	.phy_ddio_address_21(\phy_ddio_address[21] ),
	.phy_ddio_address_22(\phy_ddio_address[22] ),
	.phy_ddio_address_23(\phy_ddio_address[23] ),
	.phy_ddio_address_24(\phy_ddio_address[24] ),
	.phy_ddio_address_25(\phy_ddio_address[25] ),
	.phy_ddio_address_26(\phy_ddio_address[26] ),
	.phy_ddio_address_27(\phy_ddio_address[27] ),
	.phy_ddio_address_28(\phy_ddio_address[28] ),
	.phy_ddio_address_29(\phy_ddio_address[29] ),
	.phy_ddio_address_30(\phy_ddio_address[30] ),
	.phy_ddio_address_31(\phy_ddio_address[31] ),
	.phy_ddio_address_32(\phy_ddio_address[32] ),
	.phy_ddio_address_33(\phy_ddio_address[33] ),
	.phy_ddio_address_34(\phy_ddio_address[34] ),
	.phy_ddio_address_35(\phy_ddio_address[35] ),
	.phy_ddio_address_36(\phy_ddio_address[36] ),
	.phy_ddio_address_37(\phy_ddio_address[37] ),
	.phy_ddio_address_38(\phy_ddio_address[38] ),
	.phy_ddio_address_39(\phy_ddio_address[39] ),
	.phy_ddio_address_40(\phy_ddio_address[40] ),
	.phy_ddio_address_41(\phy_ddio_address[41] ),
	.phy_ddio_address_42(\phy_ddio_address[42] ),
	.phy_ddio_address_43(\phy_ddio_address[43] ),
	.phy_ddio_address_44(\phy_ddio_address[44] ),
	.phy_ddio_address_45(\phy_ddio_address[45] ),
	.phy_ddio_address_46(\phy_ddio_address[46] ),
	.phy_ddio_address_47(\phy_ddio_address[47] ),
	.phy_ddio_address_48(\phy_ddio_address[48] ),
	.phy_ddio_address_49(\phy_ddio_address[49] ),
	.phy_ddio_address_50(\phy_ddio_address[50] ),
	.phy_ddio_address_51(\phy_ddio_address[51] ),
	.phy_ddio_address_52(\phy_ddio_address[52] ),
	.phy_ddio_address_53(\phy_ddio_address[53] ),
	.phy_ddio_address_54(\phy_ddio_address[54] ),
	.phy_ddio_address_55(\phy_ddio_address[55] ),
	.phy_ddio_address_56(\phy_ddio_address[56] ),
	.phy_ddio_address_57(\phy_ddio_address[57] ),
	.phy_ddio_address_58(\phy_ddio_address[58] ),
	.phy_ddio_address_59(\phy_ddio_address[59] ),
	.phy_ddio_bank_0(\phy_ddio_bank[0] ),
	.phy_ddio_bank_1(\phy_ddio_bank[1] ),
	.phy_ddio_bank_2(\phy_ddio_bank[2] ),
	.phy_ddio_bank_3(\phy_ddio_bank[3] ),
	.phy_ddio_bank_4(\phy_ddio_bank[4] ),
	.phy_ddio_bank_5(\phy_ddio_bank[5] ),
	.phy_ddio_bank_6(\phy_ddio_bank[6] ),
	.phy_ddio_bank_7(\phy_ddio_bank[7] ),
	.phy_ddio_bank_8(\phy_ddio_bank[8] ),
	.phy_ddio_bank_9(\phy_ddio_bank[9] ),
	.phy_ddio_bank_10(\phy_ddio_bank[10] ),
	.phy_ddio_bank_11(\phy_ddio_bank[11] ),
	.phy_ddio_cas_n_0(\phy_ddio_cas_n[0] ),
	.phy_ddio_cas_n_1(\phy_ddio_cas_n[1] ),
	.phy_ddio_cas_n_2(\phy_ddio_cas_n[2] ),
	.phy_ddio_cas_n_3(\phy_ddio_cas_n[3] ),
	.phy_ddio_ck_0(\phy_ddio_ck[0] ),
	.phy_ddio_ck_1(\phy_ddio_ck[1] ),
	.phy_ddio_cke_0(\phy_ddio_cke[0] ),
	.phy_ddio_cke_1(\phy_ddio_cke[1] ),
	.phy_ddio_cke_2(\phy_ddio_cke[2] ),
	.phy_ddio_cke_3(\phy_ddio_cke[3] ),
	.phy_ddio_cs_n_0(\phy_ddio_cs_n[0] ),
	.phy_ddio_cs_n_1(\phy_ddio_cs_n[1] ),
	.phy_ddio_cs_n_2(\phy_ddio_cs_n[2] ),
	.phy_ddio_cs_n_3(\phy_ddio_cs_n[3] ),
	.phy_ddio_dmdout_0(\phy_ddio_dmdout[0] ),
	.phy_ddio_dmdout_1(\phy_ddio_dmdout[1] ),
	.phy_ddio_dmdout_2(\phy_ddio_dmdout[2] ),
	.phy_ddio_dmdout_3(\phy_ddio_dmdout[3] ),
	.phy_ddio_dmdout_4(\phy_ddio_dmdout[4] ),
	.phy_ddio_dmdout_5(\phy_ddio_dmdout[5] ),
	.phy_ddio_dmdout_6(\phy_ddio_dmdout[6] ),
	.phy_ddio_dmdout_7(\phy_ddio_dmdout[7] ),
	.phy_ddio_dmdout_8(\phy_ddio_dmdout[8] ),
	.phy_ddio_dmdout_9(\phy_ddio_dmdout[9] ),
	.phy_ddio_dmdout_10(\phy_ddio_dmdout[10] ),
	.phy_ddio_dmdout_11(\phy_ddio_dmdout[11] ),
	.phy_ddio_dmdout_12(\phy_ddio_dmdout[12] ),
	.phy_ddio_dmdout_13(\phy_ddio_dmdout[13] ),
	.phy_ddio_dmdout_14(\phy_ddio_dmdout[14] ),
	.phy_ddio_dmdout_15(\phy_ddio_dmdout[15] ),
	.phy_ddio_dqdout_0(\phy_ddio_dqdout[0] ),
	.phy_ddio_dqdout_1(\phy_ddio_dqdout[1] ),
	.phy_ddio_dqdout_2(\phy_ddio_dqdout[2] ),
	.phy_ddio_dqdout_3(\phy_ddio_dqdout[3] ),
	.phy_ddio_dqdout_4(\phy_ddio_dqdout[4] ),
	.phy_ddio_dqdout_5(\phy_ddio_dqdout[5] ),
	.phy_ddio_dqdout_6(\phy_ddio_dqdout[6] ),
	.phy_ddio_dqdout_7(\phy_ddio_dqdout[7] ),
	.phy_ddio_dqdout_8(\phy_ddio_dqdout[8] ),
	.phy_ddio_dqdout_9(\phy_ddio_dqdout[9] ),
	.phy_ddio_dqdout_10(\phy_ddio_dqdout[10] ),
	.phy_ddio_dqdout_11(\phy_ddio_dqdout[11] ),
	.phy_ddio_dqdout_12(\phy_ddio_dqdout[12] ),
	.phy_ddio_dqdout_13(\phy_ddio_dqdout[13] ),
	.phy_ddio_dqdout_14(\phy_ddio_dqdout[14] ),
	.phy_ddio_dqdout_15(\phy_ddio_dqdout[15] ),
	.phy_ddio_dqdout_16(\phy_ddio_dqdout[16] ),
	.phy_ddio_dqdout_17(\phy_ddio_dqdout[17] ),
	.phy_ddio_dqdout_18(\phy_ddio_dqdout[18] ),
	.phy_ddio_dqdout_19(\phy_ddio_dqdout[19] ),
	.phy_ddio_dqdout_20(\phy_ddio_dqdout[20] ),
	.phy_ddio_dqdout_21(\phy_ddio_dqdout[21] ),
	.phy_ddio_dqdout_22(\phy_ddio_dqdout[22] ),
	.phy_ddio_dqdout_23(\phy_ddio_dqdout[23] ),
	.phy_ddio_dqdout_24(\phy_ddio_dqdout[24] ),
	.phy_ddio_dqdout_25(\phy_ddio_dqdout[25] ),
	.phy_ddio_dqdout_26(\phy_ddio_dqdout[26] ),
	.phy_ddio_dqdout_27(\phy_ddio_dqdout[27] ),
	.phy_ddio_dqdout_28(\phy_ddio_dqdout[28] ),
	.phy_ddio_dqdout_29(\phy_ddio_dqdout[29] ),
	.phy_ddio_dqdout_30(\phy_ddio_dqdout[30] ),
	.phy_ddio_dqdout_31(\phy_ddio_dqdout[31] ),
	.phy_ddio_dqdout_36(\phy_ddio_dqdout[36] ),
	.phy_ddio_dqdout_37(\phy_ddio_dqdout[37] ),
	.phy_ddio_dqdout_38(\phy_ddio_dqdout[38] ),
	.phy_ddio_dqdout_39(\phy_ddio_dqdout[39] ),
	.phy_ddio_dqdout_40(\phy_ddio_dqdout[40] ),
	.phy_ddio_dqdout_41(\phy_ddio_dqdout[41] ),
	.phy_ddio_dqdout_42(\phy_ddio_dqdout[42] ),
	.phy_ddio_dqdout_43(\phy_ddio_dqdout[43] ),
	.phy_ddio_dqdout_44(\phy_ddio_dqdout[44] ),
	.phy_ddio_dqdout_45(\phy_ddio_dqdout[45] ),
	.phy_ddio_dqdout_46(\phy_ddio_dqdout[46] ),
	.phy_ddio_dqdout_47(\phy_ddio_dqdout[47] ),
	.phy_ddio_dqdout_48(\phy_ddio_dqdout[48] ),
	.phy_ddio_dqdout_49(\phy_ddio_dqdout[49] ),
	.phy_ddio_dqdout_50(\phy_ddio_dqdout[50] ),
	.phy_ddio_dqdout_51(\phy_ddio_dqdout[51] ),
	.phy_ddio_dqdout_52(\phy_ddio_dqdout[52] ),
	.phy_ddio_dqdout_53(\phy_ddio_dqdout[53] ),
	.phy_ddio_dqdout_54(\phy_ddio_dqdout[54] ),
	.phy_ddio_dqdout_55(\phy_ddio_dqdout[55] ),
	.phy_ddio_dqdout_56(\phy_ddio_dqdout[56] ),
	.phy_ddio_dqdout_57(\phy_ddio_dqdout[57] ),
	.phy_ddio_dqdout_58(\phy_ddio_dqdout[58] ),
	.phy_ddio_dqdout_59(\phy_ddio_dqdout[59] ),
	.phy_ddio_dqdout_60(\phy_ddio_dqdout[60] ),
	.phy_ddio_dqdout_61(\phy_ddio_dqdout[61] ),
	.phy_ddio_dqdout_62(\phy_ddio_dqdout[62] ),
	.phy_ddio_dqdout_63(\phy_ddio_dqdout[63] ),
	.phy_ddio_dqdout_64(\phy_ddio_dqdout[64] ),
	.phy_ddio_dqdout_65(\phy_ddio_dqdout[65] ),
	.phy_ddio_dqdout_66(\phy_ddio_dqdout[66] ),
	.phy_ddio_dqdout_67(\phy_ddio_dqdout[67] ),
	.phy_ddio_dqdout_72(\phy_ddio_dqdout[72] ),
	.phy_ddio_dqdout_73(\phy_ddio_dqdout[73] ),
	.phy_ddio_dqdout_74(\phy_ddio_dqdout[74] ),
	.phy_ddio_dqdout_75(\phy_ddio_dqdout[75] ),
	.phy_ddio_dqdout_76(\phy_ddio_dqdout[76] ),
	.phy_ddio_dqdout_77(\phy_ddio_dqdout[77] ),
	.phy_ddio_dqdout_78(\phy_ddio_dqdout[78] ),
	.phy_ddio_dqdout_79(\phy_ddio_dqdout[79] ),
	.phy_ddio_dqdout_80(\phy_ddio_dqdout[80] ),
	.phy_ddio_dqdout_81(\phy_ddio_dqdout[81] ),
	.phy_ddio_dqdout_82(\phy_ddio_dqdout[82] ),
	.phy_ddio_dqdout_83(\phy_ddio_dqdout[83] ),
	.phy_ddio_dqdout_84(\phy_ddio_dqdout[84] ),
	.phy_ddio_dqdout_85(\phy_ddio_dqdout[85] ),
	.phy_ddio_dqdout_86(\phy_ddio_dqdout[86] ),
	.phy_ddio_dqdout_87(\phy_ddio_dqdout[87] ),
	.phy_ddio_dqdout_88(\phy_ddio_dqdout[88] ),
	.phy_ddio_dqdout_89(\phy_ddio_dqdout[89] ),
	.phy_ddio_dqdout_90(\phy_ddio_dqdout[90] ),
	.phy_ddio_dqdout_91(\phy_ddio_dqdout[91] ),
	.phy_ddio_dqdout_92(\phy_ddio_dqdout[92] ),
	.phy_ddio_dqdout_93(\phy_ddio_dqdout[93] ),
	.phy_ddio_dqdout_94(\phy_ddio_dqdout[94] ),
	.phy_ddio_dqdout_95(\phy_ddio_dqdout[95] ),
	.phy_ddio_dqdout_96(\phy_ddio_dqdout[96] ),
	.phy_ddio_dqdout_97(\phy_ddio_dqdout[97] ),
	.phy_ddio_dqdout_98(\phy_ddio_dqdout[98] ),
	.phy_ddio_dqdout_99(\phy_ddio_dqdout[99] ),
	.phy_ddio_dqdout_100(\phy_ddio_dqdout[100] ),
	.phy_ddio_dqdout_101(\phy_ddio_dqdout[101] ),
	.phy_ddio_dqdout_102(\phy_ddio_dqdout[102] ),
	.phy_ddio_dqdout_103(\phy_ddio_dqdout[103] ),
	.phy_ddio_dqdout_108(\phy_ddio_dqdout[108] ),
	.phy_ddio_dqdout_109(\phy_ddio_dqdout[109] ),
	.phy_ddio_dqdout_110(\phy_ddio_dqdout[110] ),
	.phy_ddio_dqdout_111(\phy_ddio_dqdout[111] ),
	.phy_ddio_dqdout_112(\phy_ddio_dqdout[112] ),
	.phy_ddio_dqdout_113(\phy_ddio_dqdout[113] ),
	.phy_ddio_dqdout_114(\phy_ddio_dqdout[114] ),
	.phy_ddio_dqdout_115(\phy_ddio_dqdout[115] ),
	.phy_ddio_dqdout_116(\phy_ddio_dqdout[116] ),
	.phy_ddio_dqdout_117(\phy_ddio_dqdout[117] ),
	.phy_ddio_dqdout_118(\phy_ddio_dqdout[118] ),
	.phy_ddio_dqdout_119(\phy_ddio_dqdout[119] ),
	.phy_ddio_dqdout_120(\phy_ddio_dqdout[120] ),
	.phy_ddio_dqdout_121(\phy_ddio_dqdout[121] ),
	.phy_ddio_dqdout_122(\phy_ddio_dqdout[122] ),
	.phy_ddio_dqdout_123(\phy_ddio_dqdout[123] ),
	.phy_ddio_dqdout_124(\phy_ddio_dqdout[124] ),
	.phy_ddio_dqdout_125(\phy_ddio_dqdout[125] ),
	.phy_ddio_dqdout_126(\phy_ddio_dqdout[126] ),
	.phy_ddio_dqdout_127(\phy_ddio_dqdout[127] ),
	.phy_ddio_dqdout_128(\phy_ddio_dqdout[128] ),
	.phy_ddio_dqdout_129(\phy_ddio_dqdout[129] ),
	.phy_ddio_dqdout_130(\phy_ddio_dqdout[130] ),
	.phy_ddio_dqdout_131(\phy_ddio_dqdout[131] ),
	.phy_ddio_dqdout_132(\phy_ddio_dqdout[132] ),
	.phy_ddio_dqdout_133(\phy_ddio_dqdout[133] ),
	.phy_ddio_dqdout_134(\phy_ddio_dqdout[134] ),
	.phy_ddio_dqdout_135(\phy_ddio_dqdout[135] ),
	.phy_ddio_dqdout_136(\phy_ddio_dqdout[136] ),
	.phy_ddio_dqdout_137(\phy_ddio_dqdout[137] ),
	.phy_ddio_dqdout_138(\phy_ddio_dqdout[138] ),
	.phy_ddio_dqdout_139(\phy_ddio_dqdout[139] ),
	.phy_ddio_dqoe_0(\phy_ddio_dqoe[0] ),
	.phy_ddio_dqoe_1(\phy_ddio_dqoe[1] ),
	.phy_ddio_dqoe_2(\phy_ddio_dqoe[2] ),
	.phy_ddio_dqoe_3(\phy_ddio_dqoe[3] ),
	.phy_ddio_dqoe_4(\phy_ddio_dqoe[4] ),
	.phy_ddio_dqoe_5(\phy_ddio_dqoe[5] ),
	.phy_ddio_dqoe_6(\phy_ddio_dqoe[6] ),
	.phy_ddio_dqoe_7(\phy_ddio_dqoe[7] ),
	.phy_ddio_dqoe_8(\phy_ddio_dqoe[8] ),
	.phy_ddio_dqoe_9(\phy_ddio_dqoe[9] ),
	.phy_ddio_dqoe_10(\phy_ddio_dqoe[10] ),
	.phy_ddio_dqoe_11(\phy_ddio_dqoe[11] ),
	.phy_ddio_dqoe_12(\phy_ddio_dqoe[12] ),
	.phy_ddio_dqoe_13(\phy_ddio_dqoe[13] ),
	.phy_ddio_dqoe_14(\phy_ddio_dqoe[14] ),
	.phy_ddio_dqoe_15(\phy_ddio_dqoe[15] ),
	.phy_ddio_dqoe_18(\phy_ddio_dqoe[18] ),
	.phy_ddio_dqoe_19(\phy_ddio_dqoe[19] ),
	.phy_ddio_dqoe_20(\phy_ddio_dqoe[20] ),
	.phy_ddio_dqoe_21(\phy_ddio_dqoe[21] ),
	.phy_ddio_dqoe_22(\phy_ddio_dqoe[22] ),
	.phy_ddio_dqoe_23(\phy_ddio_dqoe[23] ),
	.phy_ddio_dqoe_24(\phy_ddio_dqoe[24] ),
	.phy_ddio_dqoe_25(\phy_ddio_dqoe[25] ),
	.phy_ddio_dqoe_26(\phy_ddio_dqoe[26] ),
	.phy_ddio_dqoe_27(\phy_ddio_dqoe[27] ),
	.phy_ddio_dqoe_28(\phy_ddio_dqoe[28] ),
	.phy_ddio_dqoe_29(\phy_ddio_dqoe[29] ),
	.phy_ddio_dqoe_30(\phy_ddio_dqoe[30] ),
	.phy_ddio_dqoe_31(\phy_ddio_dqoe[31] ),
	.phy_ddio_dqoe_32(\phy_ddio_dqoe[32] ),
	.phy_ddio_dqoe_33(\phy_ddio_dqoe[33] ),
	.phy_ddio_dqoe_36(\phy_ddio_dqoe[36] ),
	.phy_ddio_dqoe_37(\phy_ddio_dqoe[37] ),
	.phy_ddio_dqoe_38(\phy_ddio_dqoe[38] ),
	.phy_ddio_dqoe_39(\phy_ddio_dqoe[39] ),
	.phy_ddio_dqoe_40(\phy_ddio_dqoe[40] ),
	.phy_ddio_dqoe_41(\phy_ddio_dqoe[41] ),
	.phy_ddio_dqoe_42(\phy_ddio_dqoe[42] ),
	.phy_ddio_dqoe_43(\phy_ddio_dqoe[43] ),
	.phy_ddio_dqoe_44(\phy_ddio_dqoe[44] ),
	.phy_ddio_dqoe_45(\phy_ddio_dqoe[45] ),
	.phy_ddio_dqoe_46(\phy_ddio_dqoe[46] ),
	.phy_ddio_dqoe_47(\phy_ddio_dqoe[47] ),
	.phy_ddio_dqoe_48(\phy_ddio_dqoe[48] ),
	.phy_ddio_dqoe_49(\phy_ddio_dqoe[49] ),
	.phy_ddio_dqoe_50(\phy_ddio_dqoe[50] ),
	.phy_ddio_dqoe_51(\phy_ddio_dqoe[51] ),
	.phy_ddio_dqoe_54(\phy_ddio_dqoe[54] ),
	.phy_ddio_dqoe_55(\phy_ddio_dqoe[55] ),
	.phy_ddio_dqoe_56(\phy_ddio_dqoe[56] ),
	.phy_ddio_dqoe_57(\phy_ddio_dqoe[57] ),
	.phy_ddio_dqoe_58(\phy_ddio_dqoe[58] ),
	.phy_ddio_dqoe_59(\phy_ddio_dqoe[59] ),
	.phy_ddio_dqoe_60(\phy_ddio_dqoe[60] ),
	.phy_ddio_dqoe_61(\phy_ddio_dqoe[61] ),
	.phy_ddio_dqoe_62(\phy_ddio_dqoe[62] ),
	.phy_ddio_dqoe_63(\phy_ddio_dqoe[63] ),
	.phy_ddio_dqoe_64(\phy_ddio_dqoe[64] ),
	.phy_ddio_dqoe_65(\phy_ddio_dqoe[65] ),
	.phy_ddio_dqoe_66(\phy_ddio_dqoe[66] ),
	.phy_ddio_dqoe_67(\phy_ddio_dqoe[67] ),
	.phy_ddio_dqoe_68(\phy_ddio_dqoe[68] ),
	.phy_ddio_dqoe_69(\phy_ddio_dqoe[69] ),
	.phy_ddio_dqs_dout_0(\phy_ddio_dqs_dout[0] ),
	.phy_ddio_dqs_dout_1(\phy_ddio_dqs_dout[1] ),
	.phy_ddio_dqs_dout_2(\phy_ddio_dqs_dout[2] ),
	.phy_ddio_dqs_dout_3(\phy_ddio_dqs_dout[3] ),
	.phy_ddio_dqs_dout_4(\phy_ddio_dqs_dout[4] ),
	.phy_ddio_dqs_dout_5(\phy_ddio_dqs_dout[5] ),
	.phy_ddio_dqs_dout_6(\phy_ddio_dqs_dout[6] ),
	.phy_ddio_dqs_dout_7(\phy_ddio_dqs_dout[7] ),
	.phy_ddio_dqs_dout_8(\phy_ddio_dqs_dout[8] ),
	.phy_ddio_dqs_dout_9(\phy_ddio_dqs_dout[9] ),
	.phy_ddio_dqs_dout_10(\phy_ddio_dqs_dout[10] ),
	.phy_ddio_dqs_dout_11(\phy_ddio_dqs_dout[11] ),
	.phy_ddio_dqs_dout_12(\phy_ddio_dqs_dout[12] ),
	.phy_ddio_dqs_dout_13(\phy_ddio_dqs_dout[13] ),
	.phy_ddio_dqs_dout_14(\phy_ddio_dqs_dout[14] ),
	.phy_ddio_dqs_dout_15(\phy_ddio_dqs_dout[15] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_0(\phy_ddio_dqslogic_aclr_fifoctrl[0] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_1(\phy_ddio_dqslogic_aclr_fifoctrl[1] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_2(\phy_ddio_dqslogic_aclr_fifoctrl[2] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_3(\phy_ddio_dqslogic_aclr_fifoctrl[3] ),
	.phy_ddio_dqslogic_aclr_pstamble_0(\phy_ddio_dqslogic_aclr_pstamble[0] ),
	.phy_ddio_dqslogic_aclr_pstamble_1(\phy_ddio_dqslogic_aclr_pstamble[1] ),
	.phy_ddio_dqslogic_aclr_pstamble_2(\phy_ddio_dqslogic_aclr_pstamble[2] ),
	.phy_ddio_dqslogic_aclr_pstamble_3(\phy_ddio_dqslogic_aclr_pstamble[3] ),
	.phy_ddio_dqslogic_dqsena_0(\phy_ddio_dqslogic_dqsena[0] ),
	.phy_ddio_dqslogic_dqsena_1(\phy_ddio_dqslogic_dqsena[1] ),
	.phy_ddio_dqslogic_dqsena_2(\phy_ddio_dqslogic_dqsena[2] ),
	.phy_ddio_dqslogic_dqsena_3(\phy_ddio_dqslogic_dqsena[3] ),
	.phy_ddio_dqslogic_dqsena_4(\phy_ddio_dqslogic_dqsena[4] ),
	.phy_ddio_dqslogic_dqsena_5(\phy_ddio_dqslogic_dqsena[5] ),
	.phy_ddio_dqslogic_dqsena_6(\phy_ddio_dqslogic_dqsena[6] ),
	.phy_ddio_dqslogic_dqsena_7(\phy_ddio_dqslogic_dqsena[7] ),
	.phy_ddio_dqslogic_fiforeset_0(\phy_ddio_dqslogic_fiforeset[0] ),
	.phy_ddio_dqslogic_fiforeset_1(\phy_ddio_dqslogic_fiforeset[1] ),
	.phy_ddio_dqslogic_fiforeset_2(\phy_ddio_dqslogic_fiforeset[2] ),
	.phy_ddio_dqslogic_fiforeset_3(\phy_ddio_dqslogic_fiforeset[3] ),
	.phy_ddio_dqslogic_incrdataen_0(\phy_ddio_dqslogic_incrdataen[0] ),
	.phy_ddio_dqslogic_incrdataen_1(\phy_ddio_dqslogic_incrdataen[1] ),
	.phy_ddio_dqslogic_incrdataen_2(\phy_ddio_dqslogic_incrdataen[2] ),
	.phy_ddio_dqslogic_incrdataen_3(\phy_ddio_dqslogic_incrdataen[3] ),
	.phy_ddio_dqslogic_incrdataen_4(\phy_ddio_dqslogic_incrdataen[4] ),
	.phy_ddio_dqslogic_incrdataen_5(\phy_ddio_dqslogic_incrdataen[5] ),
	.phy_ddio_dqslogic_incrdataen_6(\phy_ddio_dqslogic_incrdataen[6] ),
	.phy_ddio_dqslogic_incrdataen_7(\phy_ddio_dqslogic_incrdataen[7] ),
	.phy_ddio_dqslogic_incwrptr_0(\phy_ddio_dqslogic_incwrptr[0] ),
	.phy_ddio_dqslogic_incwrptr_1(\phy_ddio_dqslogic_incwrptr[1] ),
	.phy_ddio_dqslogic_incwrptr_2(\phy_ddio_dqslogic_incwrptr[2] ),
	.phy_ddio_dqslogic_incwrptr_3(\phy_ddio_dqslogic_incwrptr[3] ),
	.phy_ddio_dqslogic_incwrptr_4(\phy_ddio_dqslogic_incwrptr[4] ),
	.phy_ddio_dqslogic_incwrptr_5(\phy_ddio_dqslogic_incwrptr[5] ),
	.phy_ddio_dqslogic_incwrptr_6(\phy_ddio_dqslogic_incwrptr[6] ),
	.phy_ddio_dqslogic_incwrptr_7(\phy_ddio_dqslogic_incwrptr[7] ),
	.phy_ddio_dqslogic_oct_0(\phy_ddio_dqslogic_oct[0] ),
	.phy_ddio_dqslogic_oct_1(\phy_ddio_dqslogic_oct[1] ),
	.phy_ddio_dqslogic_oct_2(\phy_ddio_dqslogic_oct[2] ),
	.phy_ddio_dqslogic_oct_3(\phy_ddio_dqslogic_oct[3] ),
	.phy_ddio_dqslogic_oct_4(\phy_ddio_dqslogic_oct[4] ),
	.phy_ddio_dqslogic_oct_5(\phy_ddio_dqslogic_oct[5] ),
	.phy_ddio_dqslogic_oct_6(\phy_ddio_dqslogic_oct[6] ),
	.phy_ddio_dqslogic_oct_7(\phy_ddio_dqslogic_oct[7] ),
	.phy_ddio_dqslogic_readlatency_0(\phy_ddio_dqslogic_readlatency[0] ),
	.phy_ddio_dqslogic_readlatency_1(\phy_ddio_dqslogic_readlatency[1] ),
	.phy_ddio_dqslogic_readlatency_2(\phy_ddio_dqslogic_readlatency[2] ),
	.phy_ddio_dqslogic_readlatency_3(\phy_ddio_dqslogic_readlatency[3] ),
	.phy_ddio_dqslogic_readlatency_4(\phy_ddio_dqslogic_readlatency[4] ),
	.phy_ddio_dqslogic_readlatency_5(\phy_ddio_dqslogic_readlatency[5] ),
	.phy_ddio_dqslogic_readlatency_6(\phy_ddio_dqslogic_readlatency[6] ),
	.phy_ddio_dqslogic_readlatency_7(\phy_ddio_dqslogic_readlatency[7] ),
	.phy_ddio_dqslogic_readlatency_8(\phy_ddio_dqslogic_readlatency[8] ),
	.phy_ddio_dqslogic_readlatency_9(\phy_ddio_dqslogic_readlatency[9] ),
	.phy_ddio_dqslogic_readlatency_10(\phy_ddio_dqslogic_readlatency[10] ),
	.phy_ddio_dqslogic_readlatency_11(\phy_ddio_dqslogic_readlatency[11] ),
	.phy_ddio_dqslogic_readlatency_12(\phy_ddio_dqslogic_readlatency[12] ),
	.phy_ddio_dqslogic_readlatency_13(\phy_ddio_dqslogic_readlatency[13] ),
	.phy_ddio_dqslogic_readlatency_14(\phy_ddio_dqslogic_readlatency[14] ),
	.phy_ddio_dqslogic_readlatency_15(\phy_ddio_dqslogic_readlatency[15] ),
	.phy_ddio_dqslogic_readlatency_16(\phy_ddio_dqslogic_readlatency[16] ),
	.phy_ddio_dqslogic_readlatency_17(\phy_ddio_dqslogic_readlatency[17] ),
	.phy_ddio_dqslogic_readlatency_18(\phy_ddio_dqslogic_readlatency[18] ),
	.phy_ddio_dqslogic_readlatency_19(\phy_ddio_dqslogic_readlatency[19] ),
	.phy_ddio_dqs_oe_0(\phy_ddio_dqs_oe[0] ),
	.phy_ddio_dqs_oe_1(\phy_ddio_dqs_oe[1] ),
	.phy_ddio_dqs_oe_2(\phy_ddio_dqs_oe[2] ),
	.phy_ddio_dqs_oe_3(\phy_ddio_dqs_oe[3] ),
	.phy_ddio_dqs_oe_4(\phy_ddio_dqs_oe[4] ),
	.phy_ddio_dqs_oe_5(\phy_ddio_dqs_oe[5] ),
	.phy_ddio_dqs_oe_6(\phy_ddio_dqs_oe[6] ),
	.phy_ddio_dqs_oe_7(\phy_ddio_dqs_oe[7] ),
	.phy_ddio_odt_0(\phy_ddio_odt[0] ),
	.phy_ddio_odt_1(\phy_ddio_odt[1] ),
	.phy_ddio_odt_2(\phy_ddio_odt[2] ),
	.phy_ddio_odt_3(\phy_ddio_odt[3] ),
	.phy_ddio_ras_n_0(\phy_ddio_ras_n[0] ),
	.phy_ddio_ras_n_1(\phy_ddio_ras_n[1] ),
	.phy_ddio_ras_n_2(\phy_ddio_ras_n[2] ),
	.phy_ddio_ras_n_3(\phy_ddio_ras_n[3] ),
	.phy_ddio_reset_n_0(\phy_ddio_reset_n[0] ),
	.phy_ddio_reset_n_1(\phy_ddio_reset_n[1] ),
	.phy_ddio_reset_n_2(\phy_ddio_reset_n[2] ),
	.phy_ddio_reset_n_3(\phy_ddio_reset_n[3] ),
	.phy_ddio_we_n_0(\phy_ddio_we_n[0] ),
	.phy_ddio_we_n_1(\phy_ddio_we_n[1] ),
	.phy_ddio_we_n_2(\phy_ddio_we_n[2] ),
	.phy_ddio_we_n_3(\phy_ddio_we_n[3] ),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.input_path_gen0read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.ddio_phy_dqslogic_rdatavalid({ddio_phy_dqslogic_rdatavalid_unconnected_wire_4,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid }),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

Computer_System_hps_sdram_p0_acv_ldc_25 memphy_ldc(
	.pll_dqs_clk(afi_clk),
	.pll_hr_clk(afi_clk),
	.afi_clk(ctl_clk),
	.avl_clk(\memphy_ldc|leveled_hr_clocks[0] ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

cyclonev_mem_phy hphy_inst(
	.aficasn(afi_cas_n[0]),
	.afimemclkdisable(afi_mem_clk_disable[0]),
	.afirasn(afi_ras_n[0]),
	.afirstn(afi_rst_n[0]),
	.afiwen(afi_we_n[0]),
	.avlread(gnd),
	.avlresetn(gnd),
	.avlwrite(gnd),
	.globalresetn(gnd),
	.iointcasnaclr(gnd),
	.iointrasnaclr(gnd),
	.iointresetnaclr(gnd),
	.iointwenaclr(gnd),
	.plladdrcmdclk(!ctl_clk),
	.pllaficlk(ctl_clk),
	.pllavlclk(\memphy_ldc|leveled_hr_clocks[0] ),
	.plllocked(gnd),
	.scanen(gnd),
	.softresetn(gnd),
	.afiaddr({afi_addr[19],afi_addr[18],afi_addr[17],afi_addr[16],afi_addr[15],afi_addr[14],afi_addr[13],afi_addr[12],afi_addr[11],afi_addr[10],afi_addr[9],afi_addr[8],afi_addr[7],afi_addr[6],afi_addr[5],afi_addr[4],afi_addr[3],afi_addr[2],afi_addr[1],afi_addr[0]}),
	.afiba({afi_ba[2],afi_ba[1],afi_ba[0]}),
	.aficke({afi_cke[1],afi_cke[0]}),
	.aficsn({afi_cs_n[1],afi_cs_n[0]}),
	.afidm({afi_dm[9],afi_dm[8],afi_dm[7],afi_dm[6],afi_dm[5],afi_dm[4],afi_dm[3],afi_dm[2],afi_dm[1],afi_dm[0]}),
	.afidqsburst({afi_dqs_burst[4],afi_dqs_burst[3],afi_dqs_burst[2],afi_dqs_burst[1],afi_dqs_burst[0]}),
	.afiodt({afi_odt[1],afi_odt[0]}),
	.afirdataen({afi_rdata_en[4],afi_rdata_en[3],afi_rdata_en[2],afi_rdata_en[1],afi_rdata_en[0]}),
	.afirdataenfull({afi_rdata_en_full[4],afi_rdata_en_full[3],afi_rdata_en_full[2],afi_rdata_en_full[1],afi_rdata_en_full[0]}),
	.afiwdata({afi_wdata[79],afi_wdata[78],afi_wdata[77],afi_wdata[76],afi_wdata[75],afi_wdata[74],afi_wdata[73],afi_wdata[72],afi_wdata[71],afi_wdata[70],afi_wdata[69],afi_wdata[68],afi_wdata[67],afi_wdata[66],afi_wdata[65],afi_wdata[64],afi_wdata[63],afi_wdata[62],afi_wdata[61],afi_wdata[60],afi_wdata[59],afi_wdata[58],afi_wdata[57],afi_wdata[56],afi_wdata[55],afi_wdata[54],afi_wdata[53],afi_wdata[52],
afi_wdata[51],afi_wdata[50],afi_wdata[49],afi_wdata[48],afi_wdata[47],afi_wdata[46],afi_wdata[45],afi_wdata[44],afi_wdata[43],afi_wdata[42],afi_wdata[41],afi_wdata[40],afi_wdata[39],afi_wdata[38],afi_wdata[37],afi_wdata[36],afi_wdata[35],afi_wdata[34],afi_wdata[33],afi_wdata[32],afi_wdata[31],afi_wdata[30],afi_wdata[29],afi_wdata[28],afi_wdata[27],afi_wdata[26],afi_wdata[25],afi_wdata[24],
afi_wdata[23],afi_wdata[22],afi_wdata[21],afi_wdata[20],afi_wdata[19],afi_wdata[18],afi_wdata[17],afi_wdata[16],afi_wdata[15],afi_wdata[14],afi_wdata[13],afi_wdata[12],afi_wdata[11],afi_wdata[10],afi_wdata[9],afi_wdata[8],afi_wdata[7],afi_wdata[6],afi_wdata[5],afi_wdata[4],afi_wdata[3],afi_wdata[2],afi_wdata[1],afi_wdata[0]}),
	.afiwdatavalid({afi_wdata_valid[4],afi_wdata_valid[3],afi_wdata_valid[2],afi_wdata_valid[1],afi_wdata_valid[0]}),
	.avladdress({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.avlwritedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfgaddlat({gnd,gnd,gnd,cfg_addlat[4],cfg_addlat[3],cfg_addlat[2],cfg_addlat[1],cfg_addlat[0]}),
	.cfgbankaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_bankaddrwidth[2],cfg_bankaddrwidth[1],cfg_bankaddrwidth[0]}),
	.cfgcaswrlat({gnd,gnd,gnd,gnd,cfg_caswrlat[3],cfg_caswrlat[2],cfg_caswrlat[1],cfg_caswrlat[0]}),
	.cfgcoladdrwidth({gnd,gnd,gnd,cfg_coladdrwidth[4],cfg_coladdrwidth[3],cfg_coladdrwidth[2],cfg_coladdrwidth[1],cfg_coladdrwidth[0]}),
	.cfgcsaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_csaddrwidth[2],cfg_csaddrwidth[1],cfg_csaddrwidth[0]}),
	.cfgdevicewidth({gnd,gnd,gnd,gnd,cfg_devicewidth[3],cfg_devicewidth[2],cfg_devicewidth[1],cfg_devicewidth[0]}),
	.cfgdramconfig({gnd,gnd,gnd,cfg_dramconfig[20],cfg_dramconfig[19],cfg_dramconfig[18],cfg_dramconfig[17],cfg_dramconfig[16],cfg_dramconfig[15],cfg_dramconfig[14],cfg_dramconfig[13],cfg_dramconfig[12],cfg_dramconfig[11],cfg_dramconfig[10],cfg_dramconfig[9],cfg_dramconfig[8],cfg_dramconfig[7],cfg_dramconfig[6],cfg_dramconfig[5],cfg_dramconfig[4],
cfg_dramconfig[3],cfg_dramconfig[2],cfg_dramconfig[1],cfg_dramconfig[0]}),
	.cfginterfacewidth({cfg_interfacewidth[7],cfg_interfacewidth[6],cfg_interfacewidth[5],cfg_interfacewidth[4],cfg_interfacewidth[3],cfg_interfacewidth[2],cfg_interfacewidth[1],cfg_interfacewidth[0]}),
	.cfgrowaddrwidth({gnd,gnd,gnd,cfg_rowaddrwidth[4],cfg_rowaddrwidth[3],cfg_rowaddrwidth[2],cfg_rowaddrwidth[1],cfg_rowaddrwidth[0]}),
	.cfgtcl({gnd,gnd,gnd,cfg_tcl[4],cfg_tcl[3],cfg_tcl[2],cfg_tcl[1],cfg_tcl[0]}),
	.cfgtmrd({gnd,gnd,gnd,gnd,cfg_tmrd[3],cfg_tmrd[2],cfg_tmrd[1],cfg_tmrd[0]}),
	.cfgtrefi({gnd,gnd,gnd,cfg_trefi[12],cfg_trefi[11],cfg_trefi[10],cfg_trefi[9],cfg_trefi[8],cfg_trefi[7],cfg_trefi[6],cfg_trefi[5],cfg_trefi[4],cfg_trefi[3],cfg_trefi[2],cfg_trefi[1],cfg_trefi[0]}),
	.cfgtrfc({cfg_trfc[7],cfg_trfc[6],cfg_trfc[5],cfg_trfc[4],cfg_trfc[3],cfg_trfc[2],cfg_trfc[1],cfg_trfc[0]}),
	.cfgtwr({gnd,gnd,gnd,gnd,cfg_twr[3],cfg_twr[2],cfg_twr[1],cfg_twr[0]}),
	.ddiophydqdin({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] }),
	.ddiophydqslogicrdatavalid({vcc,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid }),
	.iointaddraclr(16'b0000000000000000),
	.iointaddrdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointbaaclr(3'b000),
	.iointbadout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointcasndout({gnd,gnd,gnd,gnd}),
	.iointckdout({gnd,gnd,gnd,gnd}),
	.iointckeaclr(2'b00),
	.iointckedout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointckndout({gnd,gnd,gnd,gnd}),
	.iointcsnaclr(2'b00),
	.iointcsndout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdmdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqoe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iointdqsbdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsboe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicaclrfifoctrl(5'b00000),
	.iointdqslogicaclrpstamble(5'b00000),
	.iointdqslogicdqsena({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicfiforeset({gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicincrdataen({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicincwrptr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicoct({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicreadlatency({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsoe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointodtaclr(2'b00),
	.iointodtdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointrasndout({gnd,gnd,gnd,gnd}),
	.iointresetndout({gnd,gnd,gnd,gnd}),
	.iointwendout({gnd,gnd,gnd,gnd}),
	.aficalfail(afi_cal_fail),
	.aficalsuccess(afi_cal_success),
	.afirdatavalid(afi_rdata_valid[0]),
	.avlwaitrequest(),
	.ctlresetn(ctl_reset_n),
	.iointaficalfail(),
	.iointaficalsuccess(),
	.phyddiocasnaclr(),
	.phyddiorasnaclr(),
	.phyddioresetnaclr(),
	.phyddiowenaclr(),
	.phyresetn(),
	.afirdata(hphy_inst_AFIRDATA_bus),
	.afirlat(),
	.afiwlat(hphy_inst_AFIWLAT_bus),
	.avlreaddata(),
	.iointafirlat(),
	.iointafiwlat(),
	.iointdqdin(),
	.iointdqslogicrdatavalid(),
	.phyddioaddraclr(),
	.phyddioaddrdout(hphy_inst_PHYDDIOADDRDOUT_bus),
	.phyddiobaaclr(),
	.phyddiobadout(hphy_inst_PHYDDIOBADOUT_bus),
	.phyddiocasndout(hphy_inst_PHYDDIOCASNDOUT_bus),
	.phyddiockdout(hphy_inst_PHYDDIOCKDOUT_bus),
	.phyddiockeaclr(),
	.phyddiockedout(hphy_inst_PHYDDIOCKEDOUT_bus),
	.phyddiockndout(),
	.phyddiocsnaclr(),
	.phyddiocsndout(hphy_inst_PHYDDIOCSNDOUT_bus),
	.phyddiodmdout(hphy_inst_PHYDDIODMDOUT_bus),
	.phyddiodqdout(hphy_inst_PHYDDIODQDOUT_bus),
	.phyddiodqoe(hphy_inst_PHYDDIODQOE_bus),
	.phyddiodqsbdout(),
	.phyddiodqsboe(),
	.phyddiodqsdout(hphy_inst_PHYDDIODQSDOUT_bus),
	.phyddiodqslogicaclrfifoctrl(hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus),
	.phyddiodqslogicaclrpstamble(hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus),
	.phyddiodqslogicdqsena(hphy_inst_PHYDDIODQSLOGICDQSENA_bus),
	.phyddiodqslogicfiforeset(hphy_inst_PHYDDIODQSLOGICFIFORESET_bus),
	.phyddiodqslogicincrdataen(hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus),
	.phyddiodqslogicincwrptr(hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus),
	.phyddiodqslogicoct(hphy_inst_PHYDDIODQSLOGICOCT_bus),
	.phyddiodqslogicreadlatency(hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus),
	.phyddiodqsoe(hphy_inst_PHYDDIODQSOE_bus),
	.phyddioodtaclr(),
	.phyddioodtdout(hphy_inst_PHYDDIOODTDOUT_bus),
	.phyddiorasndout(hphy_inst_PHYDDIORASNDOUT_bus),
	.phyddioresetndout(hphy_inst_PHYDDIORESETNDOUT_bus),
	.phyddiowendout(hphy_inst_PHYDDIOWENDOUT_bus));
defparam hphy_inst.hphy_ac_ddr_disable = "true";
defparam hphy_inst.hphy_atpg_en = "false";
defparam hphy_inst.hphy_csr_pipelineglobalenable = "true";
defparam hphy_inst.hphy_datapath_ac_delay = "one_and_half_cycles";
defparam hphy_inst.hphy_datapath_delay = "one_cycle";
defparam hphy_inst.hphy_reset_delay_en = "false";
defparam hphy_inst.hphy_use_hphy = "true";
defparam hphy_inst.hphy_wrap_back_en = "false";
defparam hphy_inst.m_hphy_ac_rom_content = 1200'b100000011100000000000000000000100000011110000000000000000000010000000010000000010001110001010000000010000000010101110000010000000010010000000000000110010000000010100000001000011000010000000010110000000000000000010000001110000000010000000000010000000010000000010001101001010000000010000000010011101000010000000010100000000000000110010000000010010000001000011000010000000010110000000000000000110000011110000000000000000000111000011110000000000000000000110000011110000000000000000000010000011010000000000000000000010000011010110000000000000000010000001010000000010000000000010000010010000000000000000000011100100110000000000000000000011100100110110000000000000000011100100110000000000000001000011100100110110000000000001000111000111110000000000000000000111100111110000000000000000000111000011110000000000000000000011000000110000000000000000000011000100110000000000000000000010011010110000000000000000000010011010110110000000000000000010011010110000000000000001000010011010110110000000000001000110011011110000000000000000000010000010110000000000000001000010000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam hphy_inst.m_hphy_ac_rom_init_file = "hps_ac_rom.hex";
defparam hphy_inst.m_hphy_inst_rom_content = 2560'b1000000000000000000010000000011010000000000010000001100000000000100000100000000000001000001010000000000010000011000000000000100000111000000000001000000100000000000010000100100000000000100001010000000000001000010110000000000010000110000000000000100001000000000000000000100000000000000010000110100000000000000010001000000000001010011010000000100000000110100000000000000010010000000010000000011010000000000000001001100000000000101001101000000000001000011010000000100000000110100000000000000010110110100000001100110011101000000000001010111010000000100011001110100000000000101110001000000011101100100010000000000010100000100000001010110010001000100000000110100000000000110011100000000000001100110110000000000011100111000000000000000011000000000000100000110011100000001000001100111000000010000011001110000000100000110011100000000000001101000000000000000001101000000000000000011010000000000000000110100000000000000001101000000001100000111010000000011000010000100000000110000100001000000001100001000010000000000010100110100000000000100001101000000010000000011010000000000011001110000000000000110011011000000000001110011100000000000000001100000000000011000011001110000000110000110011100000001100001100111000000011000011001110000000000000110100000000000000000110100000000000000001101000000000000000011010000000000000000110100000000111000011101000000001110001000010000000011100010000100000000111000100001000000000001010011010000000000010000110100000001000000001101000000000000001000101011000000000000110110110001000000001101000000000000001000101101000000000000111111010000000000001111110100000001000011111101000010000001111111010000100000100001110100001000001000011101000010000010000111010000000000100010110100000000000011111101000000000000111111010000000101001111110100010000000011010000000010000001110100010000100000100001000100001000001000010001000010000010000100010000100000011110110100001000001000011101000010000010000111010000100000100001110100000001010011010000000010000001111111010000100000100001110100001000001000011101000010000010000111010000100000100000000100001000001000010001000010000010000100010000100000100001000100000000001000100000000000011000110100000000000100001101000000000001110011010000000100000000110100000000000000000000000000000001000000000000000000010100000000000000000110000000000000010000000000000000000000000000000100000000000100000001000000000001010000010000000000011000000100000001000000000001000000000001001000110000000000010000110100000000000101001101000000010000000011010000000010000001111000010001000000001101000000000000000000000000000;
defparam hphy_inst.m_hphy_inst_rom_init_file = "hps_inst_rom.hex";

endmodule

module Computer_System_hps_sdram_p0_acv_hard_io_pads (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	phy_ddio_address_0,
	phy_ddio_address_1,
	phy_ddio_address_2,
	phy_ddio_address_3,
	phy_ddio_address_4,
	phy_ddio_address_5,
	phy_ddio_address_6,
	phy_ddio_address_7,
	phy_ddio_address_8,
	phy_ddio_address_9,
	phy_ddio_address_10,
	phy_ddio_address_11,
	phy_ddio_address_12,
	phy_ddio_address_13,
	phy_ddio_address_14,
	phy_ddio_address_15,
	phy_ddio_address_16,
	phy_ddio_address_17,
	phy_ddio_address_18,
	phy_ddio_address_19,
	phy_ddio_address_20,
	phy_ddio_address_21,
	phy_ddio_address_22,
	phy_ddio_address_23,
	phy_ddio_address_24,
	phy_ddio_address_25,
	phy_ddio_address_26,
	phy_ddio_address_27,
	phy_ddio_address_28,
	phy_ddio_address_29,
	phy_ddio_address_30,
	phy_ddio_address_31,
	phy_ddio_address_32,
	phy_ddio_address_33,
	phy_ddio_address_34,
	phy_ddio_address_35,
	phy_ddio_address_36,
	phy_ddio_address_37,
	phy_ddio_address_38,
	phy_ddio_address_39,
	phy_ddio_address_40,
	phy_ddio_address_41,
	phy_ddio_address_42,
	phy_ddio_address_43,
	phy_ddio_address_44,
	phy_ddio_address_45,
	phy_ddio_address_46,
	phy_ddio_address_47,
	phy_ddio_address_48,
	phy_ddio_address_49,
	phy_ddio_address_50,
	phy_ddio_address_51,
	phy_ddio_address_52,
	phy_ddio_address_53,
	phy_ddio_address_54,
	phy_ddio_address_55,
	phy_ddio_address_56,
	phy_ddio_address_57,
	phy_ddio_address_58,
	phy_ddio_address_59,
	phy_ddio_bank_0,
	phy_ddio_bank_1,
	phy_ddio_bank_2,
	phy_ddio_bank_3,
	phy_ddio_bank_4,
	phy_ddio_bank_5,
	phy_ddio_bank_6,
	phy_ddio_bank_7,
	phy_ddio_bank_8,
	phy_ddio_bank_9,
	phy_ddio_bank_10,
	phy_ddio_bank_11,
	phy_ddio_cas_n_0,
	phy_ddio_cas_n_1,
	phy_ddio_cas_n_2,
	phy_ddio_cas_n_3,
	phy_ddio_ck_0,
	phy_ddio_ck_1,
	phy_ddio_cke_0,
	phy_ddio_cke_1,
	phy_ddio_cke_2,
	phy_ddio_cke_3,
	phy_ddio_cs_n_0,
	phy_ddio_cs_n_1,
	phy_ddio_cs_n_2,
	phy_ddio_cs_n_3,
	phy_ddio_dmdout_0,
	phy_ddio_dmdout_1,
	phy_ddio_dmdout_2,
	phy_ddio_dmdout_3,
	phy_ddio_dmdout_4,
	phy_ddio_dmdout_5,
	phy_ddio_dmdout_6,
	phy_ddio_dmdout_7,
	phy_ddio_dmdout_8,
	phy_ddio_dmdout_9,
	phy_ddio_dmdout_10,
	phy_ddio_dmdout_11,
	phy_ddio_dmdout_12,
	phy_ddio_dmdout_13,
	phy_ddio_dmdout_14,
	phy_ddio_dmdout_15,
	phy_ddio_dqdout_0,
	phy_ddio_dqdout_1,
	phy_ddio_dqdout_2,
	phy_ddio_dqdout_3,
	phy_ddio_dqdout_4,
	phy_ddio_dqdout_5,
	phy_ddio_dqdout_6,
	phy_ddio_dqdout_7,
	phy_ddio_dqdout_8,
	phy_ddio_dqdout_9,
	phy_ddio_dqdout_10,
	phy_ddio_dqdout_11,
	phy_ddio_dqdout_12,
	phy_ddio_dqdout_13,
	phy_ddio_dqdout_14,
	phy_ddio_dqdout_15,
	phy_ddio_dqdout_16,
	phy_ddio_dqdout_17,
	phy_ddio_dqdout_18,
	phy_ddio_dqdout_19,
	phy_ddio_dqdout_20,
	phy_ddio_dqdout_21,
	phy_ddio_dqdout_22,
	phy_ddio_dqdout_23,
	phy_ddio_dqdout_24,
	phy_ddio_dqdout_25,
	phy_ddio_dqdout_26,
	phy_ddio_dqdout_27,
	phy_ddio_dqdout_28,
	phy_ddio_dqdout_29,
	phy_ddio_dqdout_30,
	phy_ddio_dqdout_31,
	phy_ddio_dqdout_36,
	phy_ddio_dqdout_37,
	phy_ddio_dqdout_38,
	phy_ddio_dqdout_39,
	phy_ddio_dqdout_40,
	phy_ddio_dqdout_41,
	phy_ddio_dqdout_42,
	phy_ddio_dqdout_43,
	phy_ddio_dqdout_44,
	phy_ddio_dqdout_45,
	phy_ddio_dqdout_46,
	phy_ddio_dqdout_47,
	phy_ddio_dqdout_48,
	phy_ddio_dqdout_49,
	phy_ddio_dqdout_50,
	phy_ddio_dqdout_51,
	phy_ddio_dqdout_52,
	phy_ddio_dqdout_53,
	phy_ddio_dqdout_54,
	phy_ddio_dqdout_55,
	phy_ddio_dqdout_56,
	phy_ddio_dqdout_57,
	phy_ddio_dqdout_58,
	phy_ddio_dqdout_59,
	phy_ddio_dqdout_60,
	phy_ddio_dqdout_61,
	phy_ddio_dqdout_62,
	phy_ddio_dqdout_63,
	phy_ddio_dqdout_64,
	phy_ddio_dqdout_65,
	phy_ddio_dqdout_66,
	phy_ddio_dqdout_67,
	phy_ddio_dqdout_72,
	phy_ddio_dqdout_73,
	phy_ddio_dqdout_74,
	phy_ddio_dqdout_75,
	phy_ddio_dqdout_76,
	phy_ddio_dqdout_77,
	phy_ddio_dqdout_78,
	phy_ddio_dqdout_79,
	phy_ddio_dqdout_80,
	phy_ddio_dqdout_81,
	phy_ddio_dqdout_82,
	phy_ddio_dqdout_83,
	phy_ddio_dqdout_84,
	phy_ddio_dqdout_85,
	phy_ddio_dqdout_86,
	phy_ddio_dqdout_87,
	phy_ddio_dqdout_88,
	phy_ddio_dqdout_89,
	phy_ddio_dqdout_90,
	phy_ddio_dqdout_91,
	phy_ddio_dqdout_92,
	phy_ddio_dqdout_93,
	phy_ddio_dqdout_94,
	phy_ddio_dqdout_95,
	phy_ddio_dqdout_96,
	phy_ddio_dqdout_97,
	phy_ddio_dqdout_98,
	phy_ddio_dqdout_99,
	phy_ddio_dqdout_100,
	phy_ddio_dqdout_101,
	phy_ddio_dqdout_102,
	phy_ddio_dqdout_103,
	phy_ddio_dqdout_108,
	phy_ddio_dqdout_109,
	phy_ddio_dqdout_110,
	phy_ddio_dqdout_111,
	phy_ddio_dqdout_112,
	phy_ddio_dqdout_113,
	phy_ddio_dqdout_114,
	phy_ddio_dqdout_115,
	phy_ddio_dqdout_116,
	phy_ddio_dqdout_117,
	phy_ddio_dqdout_118,
	phy_ddio_dqdout_119,
	phy_ddio_dqdout_120,
	phy_ddio_dqdout_121,
	phy_ddio_dqdout_122,
	phy_ddio_dqdout_123,
	phy_ddio_dqdout_124,
	phy_ddio_dqdout_125,
	phy_ddio_dqdout_126,
	phy_ddio_dqdout_127,
	phy_ddio_dqdout_128,
	phy_ddio_dqdout_129,
	phy_ddio_dqdout_130,
	phy_ddio_dqdout_131,
	phy_ddio_dqdout_132,
	phy_ddio_dqdout_133,
	phy_ddio_dqdout_134,
	phy_ddio_dqdout_135,
	phy_ddio_dqdout_136,
	phy_ddio_dqdout_137,
	phy_ddio_dqdout_138,
	phy_ddio_dqdout_139,
	phy_ddio_dqoe_0,
	phy_ddio_dqoe_1,
	phy_ddio_dqoe_2,
	phy_ddio_dqoe_3,
	phy_ddio_dqoe_4,
	phy_ddio_dqoe_5,
	phy_ddio_dqoe_6,
	phy_ddio_dqoe_7,
	phy_ddio_dqoe_8,
	phy_ddio_dqoe_9,
	phy_ddio_dqoe_10,
	phy_ddio_dqoe_11,
	phy_ddio_dqoe_12,
	phy_ddio_dqoe_13,
	phy_ddio_dqoe_14,
	phy_ddio_dqoe_15,
	phy_ddio_dqoe_18,
	phy_ddio_dqoe_19,
	phy_ddio_dqoe_20,
	phy_ddio_dqoe_21,
	phy_ddio_dqoe_22,
	phy_ddio_dqoe_23,
	phy_ddio_dqoe_24,
	phy_ddio_dqoe_25,
	phy_ddio_dqoe_26,
	phy_ddio_dqoe_27,
	phy_ddio_dqoe_28,
	phy_ddio_dqoe_29,
	phy_ddio_dqoe_30,
	phy_ddio_dqoe_31,
	phy_ddio_dqoe_32,
	phy_ddio_dqoe_33,
	phy_ddio_dqoe_36,
	phy_ddio_dqoe_37,
	phy_ddio_dqoe_38,
	phy_ddio_dqoe_39,
	phy_ddio_dqoe_40,
	phy_ddio_dqoe_41,
	phy_ddio_dqoe_42,
	phy_ddio_dqoe_43,
	phy_ddio_dqoe_44,
	phy_ddio_dqoe_45,
	phy_ddio_dqoe_46,
	phy_ddio_dqoe_47,
	phy_ddio_dqoe_48,
	phy_ddio_dqoe_49,
	phy_ddio_dqoe_50,
	phy_ddio_dqoe_51,
	phy_ddio_dqoe_54,
	phy_ddio_dqoe_55,
	phy_ddio_dqoe_56,
	phy_ddio_dqoe_57,
	phy_ddio_dqoe_58,
	phy_ddio_dqoe_59,
	phy_ddio_dqoe_60,
	phy_ddio_dqoe_61,
	phy_ddio_dqoe_62,
	phy_ddio_dqoe_63,
	phy_ddio_dqoe_64,
	phy_ddio_dqoe_65,
	phy_ddio_dqoe_66,
	phy_ddio_dqoe_67,
	phy_ddio_dqoe_68,
	phy_ddio_dqoe_69,
	phy_ddio_dqs_dout_0,
	phy_ddio_dqs_dout_1,
	phy_ddio_dqs_dout_2,
	phy_ddio_dqs_dout_3,
	phy_ddio_dqs_dout_4,
	phy_ddio_dqs_dout_5,
	phy_ddio_dqs_dout_6,
	phy_ddio_dqs_dout_7,
	phy_ddio_dqs_dout_8,
	phy_ddio_dqs_dout_9,
	phy_ddio_dqs_dout_10,
	phy_ddio_dqs_dout_11,
	phy_ddio_dqs_dout_12,
	phy_ddio_dqs_dout_13,
	phy_ddio_dqs_dout_14,
	phy_ddio_dqs_dout_15,
	phy_ddio_dqslogic_aclr_fifoctrl_0,
	phy_ddio_dqslogic_aclr_fifoctrl_1,
	phy_ddio_dqslogic_aclr_fifoctrl_2,
	phy_ddio_dqslogic_aclr_fifoctrl_3,
	phy_ddio_dqslogic_aclr_pstamble_0,
	phy_ddio_dqslogic_aclr_pstamble_1,
	phy_ddio_dqslogic_aclr_pstamble_2,
	phy_ddio_dqslogic_aclr_pstamble_3,
	phy_ddio_dqslogic_dqsena_0,
	phy_ddio_dqslogic_dqsena_1,
	phy_ddio_dqslogic_dqsena_2,
	phy_ddio_dqslogic_dqsena_3,
	phy_ddio_dqslogic_dqsena_4,
	phy_ddio_dqslogic_dqsena_5,
	phy_ddio_dqslogic_dqsena_6,
	phy_ddio_dqslogic_dqsena_7,
	phy_ddio_dqslogic_fiforeset_0,
	phy_ddio_dqslogic_fiforeset_1,
	phy_ddio_dqslogic_fiforeset_2,
	phy_ddio_dqslogic_fiforeset_3,
	phy_ddio_dqslogic_incrdataen_0,
	phy_ddio_dqslogic_incrdataen_1,
	phy_ddio_dqslogic_incrdataen_2,
	phy_ddio_dqslogic_incrdataen_3,
	phy_ddio_dqslogic_incrdataen_4,
	phy_ddio_dqslogic_incrdataen_5,
	phy_ddio_dqslogic_incrdataen_6,
	phy_ddio_dqslogic_incrdataen_7,
	phy_ddio_dqslogic_incwrptr_0,
	phy_ddio_dqslogic_incwrptr_1,
	phy_ddio_dqslogic_incwrptr_2,
	phy_ddio_dqslogic_incwrptr_3,
	phy_ddio_dqslogic_incwrptr_4,
	phy_ddio_dqslogic_incwrptr_5,
	phy_ddio_dqslogic_incwrptr_6,
	phy_ddio_dqslogic_incwrptr_7,
	phy_ddio_dqslogic_oct_0,
	phy_ddio_dqslogic_oct_1,
	phy_ddio_dqslogic_oct_2,
	phy_ddio_dqslogic_oct_3,
	phy_ddio_dqslogic_oct_4,
	phy_ddio_dqslogic_oct_5,
	phy_ddio_dqslogic_oct_6,
	phy_ddio_dqslogic_oct_7,
	phy_ddio_dqslogic_readlatency_0,
	phy_ddio_dqslogic_readlatency_1,
	phy_ddio_dqslogic_readlatency_2,
	phy_ddio_dqslogic_readlatency_3,
	phy_ddio_dqslogic_readlatency_4,
	phy_ddio_dqslogic_readlatency_5,
	phy_ddio_dqslogic_readlatency_6,
	phy_ddio_dqslogic_readlatency_7,
	phy_ddio_dqslogic_readlatency_8,
	phy_ddio_dqslogic_readlatency_9,
	phy_ddio_dqslogic_readlatency_10,
	phy_ddio_dqslogic_readlatency_11,
	phy_ddio_dqslogic_readlatency_12,
	phy_ddio_dqslogic_readlatency_13,
	phy_ddio_dqslogic_readlatency_14,
	phy_ddio_dqslogic_readlatency_15,
	phy_ddio_dqslogic_readlatency_16,
	phy_ddio_dqslogic_readlatency_17,
	phy_ddio_dqslogic_readlatency_18,
	phy_ddio_dqslogic_readlatency_19,
	phy_ddio_dqs_oe_0,
	phy_ddio_dqs_oe_1,
	phy_ddio_dqs_oe_2,
	phy_ddio_dqs_oe_3,
	phy_ddio_dqs_oe_4,
	phy_ddio_dqs_oe_5,
	phy_ddio_dqs_oe_6,
	phy_ddio_dqs_oe_7,
	phy_ddio_odt_0,
	phy_ddio_odt_1,
	phy_ddio_odt_2,
	phy_ddio_odt_3,
	phy_ddio_ras_n_0,
	phy_ddio_ras_n_1,
	phy_ddio_ras_n_2,
	phy_ddio_ras_n_3,
	phy_ddio_reset_n_0,
	phy_ddio_reset_n_1,
	phy_ddio_reset_n_2,
	phy_ddio_reset_n_3,
	phy_ddio_we_n_0,
	phy_ddio_we_n_1,
	phy_ddio_we_n_2,
	phy_ddio_we_n_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	input_path_gen0read_fifo_out_01,
	input_path_gen0read_fifo_out_11,
	input_path_gen0read_fifo_out_21,
	input_path_gen0read_fifo_out_31,
	input_path_gen1read_fifo_out_01,
	input_path_gen1read_fifo_out_11,
	input_path_gen1read_fifo_out_21,
	input_path_gen1read_fifo_out_31,
	input_path_gen2read_fifo_out_01,
	input_path_gen2read_fifo_out_11,
	input_path_gen2read_fifo_out_21,
	input_path_gen2read_fifo_out_31,
	input_path_gen3read_fifo_out_01,
	input_path_gen3read_fifo_out_11,
	input_path_gen3read_fifo_out_21,
	input_path_gen3read_fifo_out_31,
	input_path_gen4read_fifo_out_01,
	input_path_gen4read_fifo_out_11,
	input_path_gen4read_fifo_out_21,
	input_path_gen4read_fifo_out_31,
	input_path_gen5read_fifo_out_01,
	input_path_gen5read_fifo_out_11,
	input_path_gen5read_fifo_out_21,
	input_path_gen5read_fifo_out_31,
	input_path_gen6read_fifo_out_01,
	input_path_gen6read_fifo_out_11,
	input_path_gen6read_fifo_out_21,
	input_path_gen6read_fifo_out_31,
	input_path_gen7read_fifo_out_01,
	input_path_gen7read_fifo_out_11,
	input_path_gen7read_fifo_out_21,
	input_path_gen7read_fifo_out_31,
	input_path_gen0read_fifo_out_02,
	input_path_gen0read_fifo_out_12,
	input_path_gen0read_fifo_out_22,
	input_path_gen0read_fifo_out_32,
	input_path_gen1read_fifo_out_02,
	input_path_gen1read_fifo_out_12,
	input_path_gen1read_fifo_out_22,
	input_path_gen1read_fifo_out_32,
	input_path_gen2read_fifo_out_02,
	input_path_gen2read_fifo_out_12,
	input_path_gen2read_fifo_out_22,
	input_path_gen2read_fifo_out_32,
	input_path_gen3read_fifo_out_02,
	input_path_gen3read_fifo_out_12,
	input_path_gen3read_fifo_out_22,
	input_path_gen3read_fifo_out_32,
	input_path_gen4read_fifo_out_02,
	input_path_gen4read_fifo_out_12,
	input_path_gen4read_fifo_out_22,
	input_path_gen4read_fifo_out_32,
	input_path_gen5read_fifo_out_02,
	input_path_gen5read_fifo_out_12,
	input_path_gen5read_fifo_out_22,
	input_path_gen5read_fifo_out_32,
	input_path_gen6read_fifo_out_02,
	input_path_gen6read_fifo_out_12,
	input_path_gen6read_fifo_out_22,
	input_path_gen6read_fifo_out_32,
	input_path_gen7read_fifo_out_02,
	input_path_gen7read_fifo_out_12,
	input_path_gen7read_fifo_out_22,
	input_path_gen7read_fifo_out_32,
	input_path_gen0read_fifo_out_03,
	input_path_gen0read_fifo_out_13,
	input_path_gen0read_fifo_out_23,
	input_path_gen0read_fifo_out_33,
	input_path_gen1read_fifo_out_03,
	input_path_gen1read_fifo_out_13,
	input_path_gen1read_fifo_out_23,
	input_path_gen1read_fifo_out_33,
	input_path_gen2read_fifo_out_03,
	input_path_gen2read_fifo_out_13,
	input_path_gen2read_fifo_out_23,
	input_path_gen2read_fifo_out_33,
	input_path_gen3read_fifo_out_03,
	input_path_gen3read_fifo_out_13,
	input_path_gen3read_fifo_out_23,
	input_path_gen3read_fifo_out_33,
	input_path_gen4read_fifo_out_03,
	input_path_gen4read_fifo_out_13,
	input_path_gen4read_fifo_out_23,
	input_path_gen4read_fifo_out_33,
	input_path_gen5read_fifo_out_03,
	input_path_gen5read_fifo_out_13,
	input_path_gen5read_fifo_out_23,
	input_path_gen5read_fifo_out_33,
	input_path_gen6read_fifo_out_03,
	input_path_gen6read_fifo_out_13,
	input_path_gen6read_fifo_out_23,
	input_path_gen6read_fifo_out_33,
	input_path_gen7read_fifo_out_03,
	input_path_gen7read_fifo_out_13,
	input_path_gen7read_fifo_out_23,
	input_path_gen7read_fifo_out_33,
	ddio_phy_dqslogic_rdatavalid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	phy_ddio_address_0;
input 	phy_ddio_address_1;
input 	phy_ddio_address_2;
input 	phy_ddio_address_3;
input 	phy_ddio_address_4;
input 	phy_ddio_address_5;
input 	phy_ddio_address_6;
input 	phy_ddio_address_7;
input 	phy_ddio_address_8;
input 	phy_ddio_address_9;
input 	phy_ddio_address_10;
input 	phy_ddio_address_11;
input 	phy_ddio_address_12;
input 	phy_ddio_address_13;
input 	phy_ddio_address_14;
input 	phy_ddio_address_15;
input 	phy_ddio_address_16;
input 	phy_ddio_address_17;
input 	phy_ddio_address_18;
input 	phy_ddio_address_19;
input 	phy_ddio_address_20;
input 	phy_ddio_address_21;
input 	phy_ddio_address_22;
input 	phy_ddio_address_23;
input 	phy_ddio_address_24;
input 	phy_ddio_address_25;
input 	phy_ddio_address_26;
input 	phy_ddio_address_27;
input 	phy_ddio_address_28;
input 	phy_ddio_address_29;
input 	phy_ddio_address_30;
input 	phy_ddio_address_31;
input 	phy_ddio_address_32;
input 	phy_ddio_address_33;
input 	phy_ddio_address_34;
input 	phy_ddio_address_35;
input 	phy_ddio_address_36;
input 	phy_ddio_address_37;
input 	phy_ddio_address_38;
input 	phy_ddio_address_39;
input 	phy_ddio_address_40;
input 	phy_ddio_address_41;
input 	phy_ddio_address_42;
input 	phy_ddio_address_43;
input 	phy_ddio_address_44;
input 	phy_ddio_address_45;
input 	phy_ddio_address_46;
input 	phy_ddio_address_47;
input 	phy_ddio_address_48;
input 	phy_ddio_address_49;
input 	phy_ddio_address_50;
input 	phy_ddio_address_51;
input 	phy_ddio_address_52;
input 	phy_ddio_address_53;
input 	phy_ddio_address_54;
input 	phy_ddio_address_55;
input 	phy_ddio_address_56;
input 	phy_ddio_address_57;
input 	phy_ddio_address_58;
input 	phy_ddio_address_59;
input 	phy_ddio_bank_0;
input 	phy_ddio_bank_1;
input 	phy_ddio_bank_2;
input 	phy_ddio_bank_3;
input 	phy_ddio_bank_4;
input 	phy_ddio_bank_5;
input 	phy_ddio_bank_6;
input 	phy_ddio_bank_7;
input 	phy_ddio_bank_8;
input 	phy_ddio_bank_9;
input 	phy_ddio_bank_10;
input 	phy_ddio_bank_11;
input 	phy_ddio_cas_n_0;
input 	phy_ddio_cas_n_1;
input 	phy_ddio_cas_n_2;
input 	phy_ddio_cas_n_3;
input 	phy_ddio_ck_0;
input 	phy_ddio_ck_1;
input 	phy_ddio_cke_0;
input 	phy_ddio_cke_1;
input 	phy_ddio_cke_2;
input 	phy_ddio_cke_3;
input 	phy_ddio_cs_n_0;
input 	phy_ddio_cs_n_1;
input 	phy_ddio_cs_n_2;
input 	phy_ddio_cs_n_3;
input 	phy_ddio_dmdout_0;
input 	phy_ddio_dmdout_1;
input 	phy_ddio_dmdout_2;
input 	phy_ddio_dmdout_3;
input 	phy_ddio_dmdout_4;
input 	phy_ddio_dmdout_5;
input 	phy_ddio_dmdout_6;
input 	phy_ddio_dmdout_7;
input 	phy_ddio_dmdout_8;
input 	phy_ddio_dmdout_9;
input 	phy_ddio_dmdout_10;
input 	phy_ddio_dmdout_11;
input 	phy_ddio_dmdout_12;
input 	phy_ddio_dmdout_13;
input 	phy_ddio_dmdout_14;
input 	phy_ddio_dmdout_15;
input 	phy_ddio_dqdout_0;
input 	phy_ddio_dqdout_1;
input 	phy_ddio_dqdout_2;
input 	phy_ddio_dqdout_3;
input 	phy_ddio_dqdout_4;
input 	phy_ddio_dqdout_5;
input 	phy_ddio_dqdout_6;
input 	phy_ddio_dqdout_7;
input 	phy_ddio_dqdout_8;
input 	phy_ddio_dqdout_9;
input 	phy_ddio_dqdout_10;
input 	phy_ddio_dqdout_11;
input 	phy_ddio_dqdout_12;
input 	phy_ddio_dqdout_13;
input 	phy_ddio_dqdout_14;
input 	phy_ddio_dqdout_15;
input 	phy_ddio_dqdout_16;
input 	phy_ddio_dqdout_17;
input 	phy_ddio_dqdout_18;
input 	phy_ddio_dqdout_19;
input 	phy_ddio_dqdout_20;
input 	phy_ddio_dqdout_21;
input 	phy_ddio_dqdout_22;
input 	phy_ddio_dqdout_23;
input 	phy_ddio_dqdout_24;
input 	phy_ddio_dqdout_25;
input 	phy_ddio_dqdout_26;
input 	phy_ddio_dqdout_27;
input 	phy_ddio_dqdout_28;
input 	phy_ddio_dqdout_29;
input 	phy_ddio_dqdout_30;
input 	phy_ddio_dqdout_31;
input 	phy_ddio_dqdout_36;
input 	phy_ddio_dqdout_37;
input 	phy_ddio_dqdout_38;
input 	phy_ddio_dqdout_39;
input 	phy_ddio_dqdout_40;
input 	phy_ddio_dqdout_41;
input 	phy_ddio_dqdout_42;
input 	phy_ddio_dqdout_43;
input 	phy_ddio_dqdout_44;
input 	phy_ddio_dqdout_45;
input 	phy_ddio_dqdout_46;
input 	phy_ddio_dqdout_47;
input 	phy_ddio_dqdout_48;
input 	phy_ddio_dqdout_49;
input 	phy_ddio_dqdout_50;
input 	phy_ddio_dqdout_51;
input 	phy_ddio_dqdout_52;
input 	phy_ddio_dqdout_53;
input 	phy_ddio_dqdout_54;
input 	phy_ddio_dqdout_55;
input 	phy_ddio_dqdout_56;
input 	phy_ddio_dqdout_57;
input 	phy_ddio_dqdout_58;
input 	phy_ddio_dqdout_59;
input 	phy_ddio_dqdout_60;
input 	phy_ddio_dqdout_61;
input 	phy_ddio_dqdout_62;
input 	phy_ddio_dqdout_63;
input 	phy_ddio_dqdout_64;
input 	phy_ddio_dqdout_65;
input 	phy_ddio_dqdout_66;
input 	phy_ddio_dqdout_67;
input 	phy_ddio_dqdout_72;
input 	phy_ddio_dqdout_73;
input 	phy_ddio_dqdout_74;
input 	phy_ddio_dqdout_75;
input 	phy_ddio_dqdout_76;
input 	phy_ddio_dqdout_77;
input 	phy_ddio_dqdout_78;
input 	phy_ddio_dqdout_79;
input 	phy_ddio_dqdout_80;
input 	phy_ddio_dqdout_81;
input 	phy_ddio_dqdout_82;
input 	phy_ddio_dqdout_83;
input 	phy_ddio_dqdout_84;
input 	phy_ddio_dqdout_85;
input 	phy_ddio_dqdout_86;
input 	phy_ddio_dqdout_87;
input 	phy_ddio_dqdout_88;
input 	phy_ddio_dqdout_89;
input 	phy_ddio_dqdout_90;
input 	phy_ddio_dqdout_91;
input 	phy_ddio_dqdout_92;
input 	phy_ddio_dqdout_93;
input 	phy_ddio_dqdout_94;
input 	phy_ddio_dqdout_95;
input 	phy_ddio_dqdout_96;
input 	phy_ddio_dqdout_97;
input 	phy_ddio_dqdout_98;
input 	phy_ddio_dqdout_99;
input 	phy_ddio_dqdout_100;
input 	phy_ddio_dqdout_101;
input 	phy_ddio_dqdout_102;
input 	phy_ddio_dqdout_103;
input 	phy_ddio_dqdout_108;
input 	phy_ddio_dqdout_109;
input 	phy_ddio_dqdout_110;
input 	phy_ddio_dqdout_111;
input 	phy_ddio_dqdout_112;
input 	phy_ddio_dqdout_113;
input 	phy_ddio_dqdout_114;
input 	phy_ddio_dqdout_115;
input 	phy_ddio_dqdout_116;
input 	phy_ddio_dqdout_117;
input 	phy_ddio_dqdout_118;
input 	phy_ddio_dqdout_119;
input 	phy_ddio_dqdout_120;
input 	phy_ddio_dqdout_121;
input 	phy_ddio_dqdout_122;
input 	phy_ddio_dqdout_123;
input 	phy_ddio_dqdout_124;
input 	phy_ddio_dqdout_125;
input 	phy_ddio_dqdout_126;
input 	phy_ddio_dqdout_127;
input 	phy_ddio_dqdout_128;
input 	phy_ddio_dqdout_129;
input 	phy_ddio_dqdout_130;
input 	phy_ddio_dqdout_131;
input 	phy_ddio_dqdout_132;
input 	phy_ddio_dqdout_133;
input 	phy_ddio_dqdout_134;
input 	phy_ddio_dqdout_135;
input 	phy_ddio_dqdout_136;
input 	phy_ddio_dqdout_137;
input 	phy_ddio_dqdout_138;
input 	phy_ddio_dqdout_139;
input 	phy_ddio_dqoe_0;
input 	phy_ddio_dqoe_1;
input 	phy_ddio_dqoe_2;
input 	phy_ddio_dqoe_3;
input 	phy_ddio_dqoe_4;
input 	phy_ddio_dqoe_5;
input 	phy_ddio_dqoe_6;
input 	phy_ddio_dqoe_7;
input 	phy_ddio_dqoe_8;
input 	phy_ddio_dqoe_9;
input 	phy_ddio_dqoe_10;
input 	phy_ddio_dqoe_11;
input 	phy_ddio_dqoe_12;
input 	phy_ddio_dqoe_13;
input 	phy_ddio_dqoe_14;
input 	phy_ddio_dqoe_15;
input 	phy_ddio_dqoe_18;
input 	phy_ddio_dqoe_19;
input 	phy_ddio_dqoe_20;
input 	phy_ddio_dqoe_21;
input 	phy_ddio_dqoe_22;
input 	phy_ddio_dqoe_23;
input 	phy_ddio_dqoe_24;
input 	phy_ddio_dqoe_25;
input 	phy_ddio_dqoe_26;
input 	phy_ddio_dqoe_27;
input 	phy_ddio_dqoe_28;
input 	phy_ddio_dqoe_29;
input 	phy_ddio_dqoe_30;
input 	phy_ddio_dqoe_31;
input 	phy_ddio_dqoe_32;
input 	phy_ddio_dqoe_33;
input 	phy_ddio_dqoe_36;
input 	phy_ddio_dqoe_37;
input 	phy_ddio_dqoe_38;
input 	phy_ddio_dqoe_39;
input 	phy_ddio_dqoe_40;
input 	phy_ddio_dqoe_41;
input 	phy_ddio_dqoe_42;
input 	phy_ddio_dqoe_43;
input 	phy_ddio_dqoe_44;
input 	phy_ddio_dqoe_45;
input 	phy_ddio_dqoe_46;
input 	phy_ddio_dqoe_47;
input 	phy_ddio_dqoe_48;
input 	phy_ddio_dqoe_49;
input 	phy_ddio_dqoe_50;
input 	phy_ddio_dqoe_51;
input 	phy_ddio_dqoe_54;
input 	phy_ddio_dqoe_55;
input 	phy_ddio_dqoe_56;
input 	phy_ddio_dqoe_57;
input 	phy_ddio_dqoe_58;
input 	phy_ddio_dqoe_59;
input 	phy_ddio_dqoe_60;
input 	phy_ddio_dqoe_61;
input 	phy_ddio_dqoe_62;
input 	phy_ddio_dqoe_63;
input 	phy_ddio_dqoe_64;
input 	phy_ddio_dqoe_65;
input 	phy_ddio_dqoe_66;
input 	phy_ddio_dqoe_67;
input 	phy_ddio_dqoe_68;
input 	phy_ddio_dqoe_69;
input 	phy_ddio_dqs_dout_0;
input 	phy_ddio_dqs_dout_1;
input 	phy_ddio_dqs_dout_2;
input 	phy_ddio_dqs_dout_3;
input 	phy_ddio_dqs_dout_4;
input 	phy_ddio_dqs_dout_5;
input 	phy_ddio_dqs_dout_6;
input 	phy_ddio_dqs_dout_7;
input 	phy_ddio_dqs_dout_8;
input 	phy_ddio_dqs_dout_9;
input 	phy_ddio_dqs_dout_10;
input 	phy_ddio_dqs_dout_11;
input 	phy_ddio_dqs_dout_12;
input 	phy_ddio_dqs_dout_13;
input 	phy_ddio_dqs_dout_14;
input 	phy_ddio_dqs_dout_15;
input 	phy_ddio_dqslogic_aclr_fifoctrl_0;
input 	phy_ddio_dqslogic_aclr_fifoctrl_1;
input 	phy_ddio_dqslogic_aclr_fifoctrl_2;
input 	phy_ddio_dqslogic_aclr_fifoctrl_3;
input 	phy_ddio_dqslogic_aclr_pstamble_0;
input 	phy_ddio_dqslogic_aclr_pstamble_1;
input 	phy_ddio_dqslogic_aclr_pstamble_2;
input 	phy_ddio_dqslogic_aclr_pstamble_3;
input 	phy_ddio_dqslogic_dqsena_0;
input 	phy_ddio_dqslogic_dqsena_1;
input 	phy_ddio_dqslogic_dqsena_2;
input 	phy_ddio_dqslogic_dqsena_3;
input 	phy_ddio_dqslogic_dqsena_4;
input 	phy_ddio_dqslogic_dqsena_5;
input 	phy_ddio_dqslogic_dqsena_6;
input 	phy_ddio_dqslogic_dqsena_7;
input 	phy_ddio_dqslogic_fiforeset_0;
input 	phy_ddio_dqslogic_fiforeset_1;
input 	phy_ddio_dqslogic_fiforeset_2;
input 	phy_ddio_dqslogic_fiforeset_3;
input 	phy_ddio_dqslogic_incrdataen_0;
input 	phy_ddio_dqslogic_incrdataen_1;
input 	phy_ddio_dqslogic_incrdataen_2;
input 	phy_ddio_dqslogic_incrdataen_3;
input 	phy_ddio_dqslogic_incrdataen_4;
input 	phy_ddio_dqslogic_incrdataen_5;
input 	phy_ddio_dqslogic_incrdataen_6;
input 	phy_ddio_dqslogic_incrdataen_7;
input 	phy_ddio_dqslogic_incwrptr_0;
input 	phy_ddio_dqslogic_incwrptr_1;
input 	phy_ddio_dqslogic_incwrptr_2;
input 	phy_ddio_dqslogic_incwrptr_3;
input 	phy_ddio_dqslogic_incwrptr_4;
input 	phy_ddio_dqslogic_incwrptr_5;
input 	phy_ddio_dqslogic_incwrptr_6;
input 	phy_ddio_dqslogic_incwrptr_7;
input 	phy_ddio_dqslogic_oct_0;
input 	phy_ddio_dqslogic_oct_1;
input 	phy_ddio_dqslogic_oct_2;
input 	phy_ddio_dqslogic_oct_3;
input 	phy_ddio_dqslogic_oct_4;
input 	phy_ddio_dqslogic_oct_5;
input 	phy_ddio_dqslogic_oct_6;
input 	phy_ddio_dqslogic_oct_7;
input 	phy_ddio_dqslogic_readlatency_0;
input 	phy_ddio_dqslogic_readlatency_1;
input 	phy_ddio_dqslogic_readlatency_2;
input 	phy_ddio_dqslogic_readlatency_3;
input 	phy_ddio_dqslogic_readlatency_4;
input 	phy_ddio_dqslogic_readlatency_5;
input 	phy_ddio_dqslogic_readlatency_6;
input 	phy_ddio_dqslogic_readlatency_7;
input 	phy_ddio_dqslogic_readlatency_8;
input 	phy_ddio_dqslogic_readlatency_9;
input 	phy_ddio_dqslogic_readlatency_10;
input 	phy_ddio_dqslogic_readlatency_11;
input 	phy_ddio_dqslogic_readlatency_12;
input 	phy_ddio_dqslogic_readlatency_13;
input 	phy_ddio_dqslogic_readlatency_14;
input 	phy_ddio_dqslogic_readlatency_15;
input 	phy_ddio_dqslogic_readlatency_16;
input 	phy_ddio_dqslogic_readlatency_17;
input 	phy_ddio_dqslogic_readlatency_18;
input 	phy_ddio_dqslogic_readlatency_19;
input 	phy_ddio_dqs_oe_0;
input 	phy_ddio_dqs_oe_1;
input 	phy_ddio_dqs_oe_2;
input 	phy_ddio_dqs_oe_3;
input 	phy_ddio_dqs_oe_4;
input 	phy_ddio_dqs_oe_5;
input 	phy_ddio_dqs_oe_6;
input 	phy_ddio_dqs_oe_7;
input 	phy_ddio_odt_0;
input 	phy_ddio_odt_1;
input 	phy_ddio_odt_2;
input 	phy_ddio_odt_3;
input 	phy_ddio_ras_n_0;
input 	phy_ddio_ras_n_1;
input 	phy_ddio_ras_n_2;
input 	phy_ddio_ras_n_3;
input 	phy_ddio_reset_n_0;
input 	phy_ddio_reset_n_1;
input 	phy_ddio_reset_n_2;
input 	phy_ddio_reset_n_3;
input 	phy_ddio_we_n_0;
input 	phy_ddio_we_n_1;
input 	phy_ddio_we_n_2;
input 	phy_ddio_we_n_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	input_path_gen0read_fifo_out_01;
output 	input_path_gen0read_fifo_out_11;
output 	input_path_gen0read_fifo_out_21;
output 	input_path_gen0read_fifo_out_31;
output 	input_path_gen1read_fifo_out_01;
output 	input_path_gen1read_fifo_out_11;
output 	input_path_gen1read_fifo_out_21;
output 	input_path_gen1read_fifo_out_31;
output 	input_path_gen2read_fifo_out_01;
output 	input_path_gen2read_fifo_out_11;
output 	input_path_gen2read_fifo_out_21;
output 	input_path_gen2read_fifo_out_31;
output 	input_path_gen3read_fifo_out_01;
output 	input_path_gen3read_fifo_out_11;
output 	input_path_gen3read_fifo_out_21;
output 	input_path_gen3read_fifo_out_31;
output 	input_path_gen4read_fifo_out_01;
output 	input_path_gen4read_fifo_out_11;
output 	input_path_gen4read_fifo_out_21;
output 	input_path_gen4read_fifo_out_31;
output 	input_path_gen5read_fifo_out_01;
output 	input_path_gen5read_fifo_out_11;
output 	input_path_gen5read_fifo_out_21;
output 	input_path_gen5read_fifo_out_31;
output 	input_path_gen6read_fifo_out_01;
output 	input_path_gen6read_fifo_out_11;
output 	input_path_gen6read_fifo_out_21;
output 	input_path_gen6read_fifo_out_31;
output 	input_path_gen7read_fifo_out_01;
output 	input_path_gen7read_fifo_out_11;
output 	input_path_gen7read_fifo_out_21;
output 	input_path_gen7read_fifo_out_31;
output 	input_path_gen0read_fifo_out_02;
output 	input_path_gen0read_fifo_out_12;
output 	input_path_gen0read_fifo_out_22;
output 	input_path_gen0read_fifo_out_32;
output 	input_path_gen1read_fifo_out_02;
output 	input_path_gen1read_fifo_out_12;
output 	input_path_gen1read_fifo_out_22;
output 	input_path_gen1read_fifo_out_32;
output 	input_path_gen2read_fifo_out_02;
output 	input_path_gen2read_fifo_out_12;
output 	input_path_gen2read_fifo_out_22;
output 	input_path_gen2read_fifo_out_32;
output 	input_path_gen3read_fifo_out_02;
output 	input_path_gen3read_fifo_out_12;
output 	input_path_gen3read_fifo_out_22;
output 	input_path_gen3read_fifo_out_32;
output 	input_path_gen4read_fifo_out_02;
output 	input_path_gen4read_fifo_out_12;
output 	input_path_gen4read_fifo_out_22;
output 	input_path_gen4read_fifo_out_32;
output 	input_path_gen5read_fifo_out_02;
output 	input_path_gen5read_fifo_out_12;
output 	input_path_gen5read_fifo_out_22;
output 	input_path_gen5read_fifo_out_32;
output 	input_path_gen6read_fifo_out_02;
output 	input_path_gen6read_fifo_out_12;
output 	input_path_gen6read_fifo_out_22;
output 	input_path_gen6read_fifo_out_32;
output 	input_path_gen7read_fifo_out_02;
output 	input_path_gen7read_fifo_out_12;
output 	input_path_gen7read_fifo_out_22;
output 	input_path_gen7read_fifo_out_32;
output 	input_path_gen0read_fifo_out_03;
output 	input_path_gen0read_fifo_out_13;
output 	input_path_gen0read_fifo_out_23;
output 	input_path_gen0read_fifo_out_33;
output 	input_path_gen1read_fifo_out_03;
output 	input_path_gen1read_fifo_out_13;
output 	input_path_gen1read_fifo_out_23;
output 	input_path_gen1read_fifo_out_33;
output 	input_path_gen2read_fifo_out_03;
output 	input_path_gen2read_fifo_out_13;
output 	input_path_gen2read_fifo_out_23;
output 	input_path_gen2read_fifo_out_33;
output 	input_path_gen3read_fifo_out_03;
output 	input_path_gen3read_fifo_out_13;
output 	input_path_gen3read_fifo_out_23;
output 	input_path_gen3read_fifo_out_33;
output 	input_path_gen4read_fifo_out_03;
output 	input_path_gen4read_fifo_out_13;
output 	input_path_gen4read_fifo_out_23;
output 	input_path_gen4read_fifo_out_33;
output 	input_path_gen5read_fifo_out_03;
output 	input_path_gen5read_fifo_out_13;
output 	input_path_gen5read_fifo_out_23;
output 	input_path_gen5read_fifo_out_33;
output 	input_path_gen6read_fifo_out_03;
output 	input_path_gen6read_fifo_out_13;
output 	input_path_gen6read_fifo_out_23;
output 	input_path_gen6read_fifo_out_33;
output 	input_path_gen7read_fifo_out_03;
output 	input_path_gen7read_fifo_out_13;
output 	input_path_gen7read_fifo_out_23;
output 	input_path_gen7read_fifo_out_33;
output 	[4:0] ddio_phy_dqslogic_rdatavalid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_hps_sdram_p0_altdqdqs_3 \dq_ddio[3].ubidir_dq_dqs (
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.phy_ddio_dmdout_12(phy_ddio_dmdout_12),
	.phy_ddio_dmdout_13(phy_ddio_dmdout_13),
	.phy_ddio_dmdout_14(phy_ddio_dmdout_14),
	.phy_ddio_dmdout_15(phy_ddio_dmdout_15),
	.phy_ddio_dqdout_108(phy_ddio_dqdout_108),
	.phy_ddio_dqdout_109(phy_ddio_dqdout_109),
	.phy_ddio_dqdout_110(phy_ddio_dqdout_110),
	.phy_ddio_dqdout_111(phy_ddio_dqdout_111),
	.phy_ddio_dqdout_112(phy_ddio_dqdout_112),
	.phy_ddio_dqdout_113(phy_ddio_dqdout_113),
	.phy_ddio_dqdout_114(phy_ddio_dqdout_114),
	.phy_ddio_dqdout_115(phy_ddio_dqdout_115),
	.phy_ddio_dqdout_116(phy_ddio_dqdout_116),
	.phy_ddio_dqdout_117(phy_ddio_dqdout_117),
	.phy_ddio_dqdout_118(phy_ddio_dqdout_118),
	.phy_ddio_dqdout_119(phy_ddio_dqdout_119),
	.phy_ddio_dqdout_120(phy_ddio_dqdout_120),
	.phy_ddio_dqdout_121(phy_ddio_dqdout_121),
	.phy_ddio_dqdout_122(phy_ddio_dqdout_122),
	.phy_ddio_dqdout_123(phy_ddio_dqdout_123),
	.phy_ddio_dqdout_124(phy_ddio_dqdout_124),
	.phy_ddio_dqdout_125(phy_ddio_dqdout_125),
	.phy_ddio_dqdout_126(phy_ddio_dqdout_126),
	.phy_ddio_dqdout_127(phy_ddio_dqdout_127),
	.phy_ddio_dqdout_128(phy_ddio_dqdout_128),
	.phy_ddio_dqdout_129(phy_ddio_dqdout_129),
	.phy_ddio_dqdout_130(phy_ddio_dqdout_130),
	.phy_ddio_dqdout_131(phy_ddio_dqdout_131),
	.phy_ddio_dqdout_132(phy_ddio_dqdout_132),
	.phy_ddio_dqdout_133(phy_ddio_dqdout_133),
	.phy_ddio_dqdout_134(phy_ddio_dqdout_134),
	.phy_ddio_dqdout_135(phy_ddio_dqdout_135),
	.phy_ddio_dqdout_136(phy_ddio_dqdout_136),
	.phy_ddio_dqdout_137(phy_ddio_dqdout_137),
	.phy_ddio_dqdout_138(phy_ddio_dqdout_138),
	.phy_ddio_dqdout_139(phy_ddio_dqdout_139),
	.phy_ddio_dqoe_54(phy_ddio_dqoe_54),
	.phy_ddio_dqoe_55(phy_ddio_dqoe_55),
	.phy_ddio_dqoe_56(phy_ddio_dqoe_56),
	.phy_ddio_dqoe_57(phy_ddio_dqoe_57),
	.phy_ddio_dqoe_58(phy_ddio_dqoe_58),
	.phy_ddio_dqoe_59(phy_ddio_dqoe_59),
	.phy_ddio_dqoe_60(phy_ddio_dqoe_60),
	.phy_ddio_dqoe_61(phy_ddio_dqoe_61),
	.phy_ddio_dqoe_62(phy_ddio_dqoe_62),
	.phy_ddio_dqoe_63(phy_ddio_dqoe_63),
	.phy_ddio_dqoe_64(phy_ddio_dqoe_64),
	.phy_ddio_dqoe_65(phy_ddio_dqoe_65),
	.phy_ddio_dqoe_66(phy_ddio_dqoe_66),
	.phy_ddio_dqoe_67(phy_ddio_dqoe_67),
	.phy_ddio_dqoe_68(phy_ddio_dqoe_68),
	.phy_ddio_dqoe_69(phy_ddio_dqoe_69),
	.phy_ddio_dqs_dout_12(phy_ddio_dqs_dout_12),
	.phy_ddio_dqs_dout_13(phy_ddio_dqs_dout_13),
	.phy_ddio_dqs_dout_14(phy_ddio_dqs_dout_14),
	.phy_ddio_dqs_dout_15(phy_ddio_dqs_dout_15),
	.phy_ddio_dqslogic_aclr_fifoctrl_3(phy_ddio_dqslogic_aclr_fifoctrl_3),
	.phy_ddio_dqslogic_aclr_pstamble_3(phy_ddio_dqslogic_aclr_pstamble_3),
	.phy_ddio_dqslogic_dqsena_6(phy_ddio_dqslogic_dqsena_6),
	.phy_ddio_dqslogic_dqsena_7(phy_ddio_dqslogic_dqsena_7),
	.phy_ddio_dqslogic_fiforeset_3(phy_ddio_dqslogic_fiforeset_3),
	.phy_ddio_dqslogic_incrdataen_6(phy_ddio_dqslogic_incrdataen_6),
	.phy_ddio_dqslogic_incrdataen_7(phy_ddio_dqslogic_incrdataen_7),
	.phy_ddio_dqslogic_incwrptr_6(phy_ddio_dqslogic_incwrptr_6),
	.phy_ddio_dqslogic_incwrptr_7(phy_ddio_dqslogic_incwrptr_7),
	.phy_ddio_dqslogic_oct_6(phy_ddio_dqslogic_oct_6),
	.phy_ddio_dqslogic_oct_7(phy_ddio_dqslogic_oct_7),
	.phy_ddio_dqslogic_readlatency_15(phy_ddio_dqslogic_readlatency_15),
	.phy_ddio_dqslogic_readlatency_16(phy_ddio_dqslogic_readlatency_16),
	.phy_ddio_dqslogic_readlatency_17(phy_ddio_dqslogic_readlatency_17),
	.phy_ddio_dqslogic_readlatency_18(phy_ddio_dqslogic_readlatency_18),
	.phy_ddio_dqslogic_readlatency_19(phy_ddio_dqslogic_readlatency_19),
	.phy_ddio_dqs_oe_6(phy_ddio_dqs_oe_6),
	.phy_ddio_dqs_oe_7(phy_ddio_dqs_oe_7),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_13),
	.delayed_oct(delayed_oct3),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_13),
	.os(os3),
	.os_bar(os_bar3),
	.diff_oe(diff_oe3),
	.diff_oe_bar(diff_oe_bar3),
	.diff_dtc(diff_dtc3),
	.diff_dtc_bar(diff_dtc_bar3),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_03),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_13),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_23),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_33),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_03),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_13),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_23),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_33),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_03),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_13),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_23),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_33),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_03),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_13),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_23),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_33),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_03),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_13),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_23),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_33),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_03),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_13),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_23),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_33),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_03),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_13),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_23),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_33),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_03),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_13),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_23),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_33),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[3]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

Computer_System_hps_sdram_p0_altdqdqs_2 \dq_ddio[2].ubidir_dq_dqs (
	.dqsin(dqsin1),
	.pad_gen0raw_input(pad_gen0raw_input1),
	.pad_gen1raw_input(pad_gen1raw_input1),
	.pad_gen2raw_input(pad_gen2raw_input1),
	.pad_gen3raw_input(pad_gen3raw_input1),
	.pad_gen4raw_input(pad_gen4raw_input1),
	.pad_gen5raw_input(pad_gen5raw_input1),
	.pad_gen6raw_input(pad_gen6raw_input1),
	.pad_gen7raw_input(pad_gen7raw_input1),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out1),
	.phy_ddio_dmdout_8(phy_ddio_dmdout_8),
	.phy_ddio_dmdout_9(phy_ddio_dmdout_9),
	.phy_ddio_dmdout_10(phy_ddio_dmdout_10),
	.phy_ddio_dmdout_11(phy_ddio_dmdout_11),
	.phy_ddio_dqdout_72(phy_ddio_dqdout_72),
	.phy_ddio_dqdout_73(phy_ddio_dqdout_73),
	.phy_ddio_dqdout_74(phy_ddio_dqdout_74),
	.phy_ddio_dqdout_75(phy_ddio_dqdout_75),
	.phy_ddio_dqdout_76(phy_ddio_dqdout_76),
	.phy_ddio_dqdout_77(phy_ddio_dqdout_77),
	.phy_ddio_dqdout_78(phy_ddio_dqdout_78),
	.phy_ddio_dqdout_79(phy_ddio_dqdout_79),
	.phy_ddio_dqdout_80(phy_ddio_dqdout_80),
	.phy_ddio_dqdout_81(phy_ddio_dqdout_81),
	.phy_ddio_dqdout_82(phy_ddio_dqdout_82),
	.phy_ddio_dqdout_83(phy_ddio_dqdout_83),
	.phy_ddio_dqdout_84(phy_ddio_dqdout_84),
	.phy_ddio_dqdout_85(phy_ddio_dqdout_85),
	.phy_ddio_dqdout_86(phy_ddio_dqdout_86),
	.phy_ddio_dqdout_87(phy_ddio_dqdout_87),
	.phy_ddio_dqdout_88(phy_ddio_dqdout_88),
	.phy_ddio_dqdout_89(phy_ddio_dqdout_89),
	.phy_ddio_dqdout_90(phy_ddio_dqdout_90),
	.phy_ddio_dqdout_91(phy_ddio_dqdout_91),
	.phy_ddio_dqdout_92(phy_ddio_dqdout_92),
	.phy_ddio_dqdout_93(phy_ddio_dqdout_93),
	.phy_ddio_dqdout_94(phy_ddio_dqdout_94),
	.phy_ddio_dqdout_95(phy_ddio_dqdout_95),
	.phy_ddio_dqdout_96(phy_ddio_dqdout_96),
	.phy_ddio_dqdout_97(phy_ddio_dqdout_97),
	.phy_ddio_dqdout_98(phy_ddio_dqdout_98),
	.phy_ddio_dqdout_99(phy_ddio_dqdout_99),
	.phy_ddio_dqdout_100(phy_ddio_dqdout_100),
	.phy_ddio_dqdout_101(phy_ddio_dqdout_101),
	.phy_ddio_dqdout_102(phy_ddio_dqdout_102),
	.phy_ddio_dqdout_103(phy_ddio_dqdout_103),
	.phy_ddio_dqoe_36(phy_ddio_dqoe_36),
	.phy_ddio_dqoe_37(phy_ddio_dqoe_37),
	.phy_ddio_dqoe_38(phy_ddio_dqoe_38),
	.phy_ddio_dqoe_39(phy_ddio_dqoe_39),
	.phy_ddio_dqoe_40(phy_ddio_dqoe_40),
	.phy_ddio_dqoe_41(phy_ddio_dqoe_41),
	.phy_ddio_dqoe_42(phy_ddio_dqoe_42),
	.phy_ddio_dqoe_43(phy_ddio_dqoe_43),
	.phy_ddio_dqoe_44(phy_ddio_dqoe_44),
	.phy_ddio_dqoe_45(phy_ddio_dqoe_45),
	.phy_ddio_dqoe_46(phy_ddio_dqoe_46),
	.phy_ddio_dqoe_47(phy_ddio_dqoe_47),
	.phy_ddio_dqoe_48(phy_ddio_dqoe_48),
	.phy_ddio_dqoe_49(phy_ddio_dqoe_49),
	.phy_ddio_dqoe_50(phy_ddio_dqoe_50),
	.phy_ddio_dqoe_51(phy_ddio_dqoe_51),
	.phy_ddio_dqs_dout_8(phy_ddio_dqs_dout_8),
	.phy_ddio_dqs_dout_9(phy_ddio_dqs_dout_9),
	.phy_ddio_dqs_dout_10(phy_ddio_dqs_dout_10),
	.phy_ddio_dqs_dout_11(phy_ddio_dqs_dout_11),
	.phy_ddio_dqslogic_aclr_fifoctrl_2(phy_ddio_dqslogic_aclr_fifoctrl_2),
	.phy_ddio_dqslogic_aclr_pstamble_2(phy_ddio_dqslogic_aclr_pstamble_2),
	.phy_ddio_dqslogic_dqsena_4(phy_ddio_dqslogic_dqsena_4),
	.phy_ddio_dqslogic_dqsena_5(phy_ddio_dqslogic_dqsena_5),
	.phy_ddio_dqslogic_fiforeset_2(phy_ddio_dqslogic_fiforeset_2),
	.phy_ddio_dqslogic_incrdataen_4(phy_ddio_dqslogic_incrdataen_4),
	.phy_ddio_dqslogic_incrdataen_5(phy_ddio_dqslogic_incrdataen_5),
	.phy_ddio_dqslogic_incwrptr_4(phy_ddio_dqslogic_incwrptr_4),
	.phy_ddio_dqslogic_incwrptr_5(phy_ddio_dqslogic_incwrptr_5),
	.phy_ddio_dqslogic_oct_4(phy_ddio_dqslogic_oct_4),
	.phy_ddio_dqslogic_oct_5(phy_ddio_dqslogic_oct_5),
	.phy_ddio_dqslogic_readlatency_10(phy_ddio_dqslogic_readlatency_10),
	.phy_ddio_dqslogic_readlatency_11(phy_ddio_dqslogic_readlatency_11),
	.phy_ddio_dqslogic_readlatency_12(phy_ddio_dqslogic_readlatency_12),
	.phy_ddio_dqslogic_readlatency_13(phy_ddio_dqslogic_readlatency_13),
	.phy_ddio_dqslogic_readlatency_14(phy_ddio_dqslogic_readlatency_14),
	.phy_ddio_dqs_oe_4(phy_ddio_dqs_oe_4),
	.phy_ddio_dqs_oe_5(phy_ddio_dqs_oe_5),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_12),
	.delayed_oct(delayed_oct2),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_12),
	.os(os2),
	.os_bar(os_bar2),
	.diff_oe(diff_oe2),
	.diff_oe_bar(diff_oe_bar2),
	.diff_dtc(diff_dtc2),
	.diff_dtc_bar(diff_dtc_bar2),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_02),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_12),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_22),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_32),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_02),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_12),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_22),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_32),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_02),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_12),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_22),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_32),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_02),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_12),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_22),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_32),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_02),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_12),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_22),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_32),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_02),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_12),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_22),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_32),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_02),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_12),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_22),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_32),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_02),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_12),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_22),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_32),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[2]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

Computer_System_hps_sdram_p0_altdqdqs_1 \dq_ddio[1].ubidir_dq_dqs (
	.dqsin(dqsin2),
	.pad_gen0raw_input(pad_gen0raw_input2),
	.pad_gen1raw_input(pad_gen1raw_input2),
	.pad_gen2raw_input(pad_gen2raw_input2),
	.pad_gen3raw_input(pad_gen3raw_input2),
	.pad_gen4raw_input(pad_gen4raw_input2),
	.pad_gen5raw_input(pad_gen5raw_input2),
	.pad_gen6raw_input(pad_gen6raw_input2),
	.pad_gen7raw_input(pad_gen7raw_input2),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out2),
	.phy_ddio_dmdout_4(phy_ddio_dmdout_4),
	.phy_ddio_dmdout_5(phy_ddio_dmdout_5),
	.phy_ddio_dmdout_6(phy_ddio_dmdout_6),
	.phy_ddio_dmdout_7(phy_ddio_dmdout_7),
	.phy_ddio_dqdout_36(phy_ddio_dqdout_36),
	.phy_ddio_dqdout_37(phy_ddio_dqdout_37),
	.phy_ddio_dqdout_38(phy_ddio_dqdout_38),
	.phy_ddio_dqdout_39(phy_ddio_dqdout_39),
	.phy_ddio_dqdout_40(phy_ddio_dqdout_40),
	.phy_ddio_dqdout_41(phy_ddio_dqdout_41),
	.phy_ddio_dqdout_42(phy_ddio_dqdout_42),
	.phy_ddio_dqdout_43(phy_ddio_dqdout_43),
	.phy_ddio_dqdout_44(phy_ddio_dqdout_44),
	.phy_ddio_dqdout_45(phy_ddio_dqdout_45),
	.phy_ddio_dqdout_46(phy_ddio_dqdout_46),
	.phy_ddio_dqdout_47(phy_ddio_dqdout_47),
	.phy_ddio_dqdout_48(phy_ddio_dqdout_48),
	.phy_ddio_dqdout_49(phy_ddio_dqdout_49),
	.phy_ddio_dqdout_50(phy_ddio_dqdout_50),
	.phy_ddio_dqdout_51(phy_ddio_dqdout_51),
	.phy_ddio_dqdout_52(phy_ddio_dqdout_52),
	.phy_ddio_dqdout_53(phy_ddio_dqdout_53),
	.phy_ddio_dqdout_54(phy_ddio_dqdout_54),
	.phy_ddio_dqdout_55(phy_ddio_dqdout_55),
	.phy_ddio_dqdout_56(phy_ddio_dqdout_56),
	.phy_ddio_dqdout_57(phy_ddio_dqdout_57),
	.phy_ddio_dqdout_58(phy_ddio_dqdout_58),
	.phy_ddio_dqdout_59(phy_ddio_dqdout_59),
	.phy_ddio_dqdout_60(phy_ddio_dqdout_60),
	.phy_ddio_dqdout_61(phy_ddio_dqdout_61),
	.phy_ddio_dqdout_62(phy_ddio_dqdout_62),
	.phy_ddio_dqdout_63(phy_ddio_dqdout_63),
	.phy_ddio_dqdout_64(phy_ddio_dqdout_64),
	.phy_ddio_dqdout_65(phy_ddio_dqdout_65),
	.phy_ddio_dqdout_66(phy_ddio_dqdout_66),
	.phy_ddio_dqdout_67(phy_ddio_dqdout_67),
	.phy_ddio_dqoe_18(phy_ddio_dqoe_18),
	.phy_ddio_dqoe_19(phy_ddio_dqoe_19),
	.phy_ddio_dqoe_20(phy_ddio_dqoe_20),
	.phy_ddio_dqoe_21(phy_ddio_dqoe_21),
	.phy_ddio_dqoe_22(phy_ddio_dqoe_22),
	.phy_ddio_dqoe_23(phy_ddio_dqoe_23),
	.phy_ddio_dqoe_24(phy_ddio_dqoe_24),
	.phy_ddio_dqoe_25(phy_ddio_dqoe_25),
	.phy_ddio_dqoe_26(phy_ddio_dqoe_26),
	.phy_ddio_dqoe_27(phy_ddio_dqoe_27),
	.phy_ddio_dqoe_28(phy_ddio_dqoe_28),
	.phy_ddio_dqoe_29(phy_ddio_dqoe_29),
	.phy_ddio_dqoe_30(phy_ddio_dqoe_30),
	.phy_ddio_dqoe_31(phy_ddio_dqoe_31),
	.phy_ddio_dqoe_32(phy_ddio_dqoe_32),
	.phy_ddio_dqoe_33(phy_ddio_dqoe_33),
	.phy_ddio_dqs_dout_4(phy_ddio_dqs_dout_4),
	.phy_ddio_dqs_dout_5(phy_ddio_dqs_dout_5),
	.phy_ddio_dqs_dout_6(phy_ddio_dqs_dout_6),
	.phy_ddio_dqs_dout_7(phy_ddio_dqs_dout_7),
	.phy_ddio_dqslogic_aclr_fifoctrl_1(phy_ddio_dqslogic_aclr_fifoctrl_1),
	.phy_ddio_dqslogic_aclr_pstamble_1(phy_ddio_dqslogic_aclr_pstamble_1),
	.phy_ddio_dqslogic_dqsena_2(phy_ddio_dqslogic_dqsena_2),
	.phy_ddio_dqslogic_dqsena_3(phy_ddio_dqslogic_dqsena_3),
	.phy_ddio_dqslogic_fiforeset_1(phy_ddio_dqslogic_fiforeset_1),
	.phy_ddio_dqslogic_incrdataen_2(phy_ddio_dqslogic_incrdataen_2),
	.phy_ddio_dqslogic_incrdataen_3(phy_ddio_dqslogic_incrdataen_3),
	.phy_ddio_dqslogic_incwrptr_2(phy_ddio_dqslogic_incwrptr_2),
	.phy_ddio_dqslogic_incwrptr_3(phy_ddio_dqslogic_incwrptr_3),
	.phy_ddio_dqslogic_oct_2(phy_ddio_dqslogic_oct_2),
	.phy_ddio_dqslogic_oct_3(phy_ddio_dqslogic_oct_3),
	.phy_ddio_dqslogic_readlatency_5(phy_ddio_dqslogic_readlatency_5),
	.phy_ddio_dqslogic_readlatency_6(phy_ddio_dqslogic_readlatency_6),
	.phy_ddio_dqslogic_readlatency_7(phy_ddio_dqslogic_readlatency_7),
	.phy_ddio_dqslogic_readlatency_8(phy_ddio_dqslogic_readlatency_8),
	.phy_ddio_dqslogic_readlatency_9(phy_ddio_dqslogic_readlatency_9),
	.phy_ddio_dqs_oe_2(phy_ddio_dqs_oe_2),
	.phy_ddio_dqs_oe_3(phy_ddio_dqs_oe_3),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_11),
	.delayed_oct(delayed_oct1),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_11),
	.os(os1),
	.os_bar(os_bar1),
	.diff_oe(diff_oe1),
	.diff_oe_bar(diff_oe_bar1),
	.diff_dtc(diff_dtc1),
	.diff_dtc_bar(diff_dtc_bar1),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_01),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_11),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_21),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_31),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_01),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_11),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_21),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_31),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_01),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_11),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_21),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_31),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_01),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_11),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_21),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_31),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_01),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_11),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_21),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_31),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_01),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_11),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_21),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_31),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_01),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_11),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_21),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_31),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_01),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_11),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_21),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_31),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[1]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

Computer_System_hps_sdram_p0_altdqdqs \dq_ddio[0].ubidir_dq_dqs (
	.dqsin(dqsin3),
	.pad_gen0raw_input(pad_gen0raw_input3),
	.pad_gen1raw_input(pad_gen1raw_input3),
	.pad_gen2raw_input(pad_gen2raw_input3),
	.pad_gen3raw_input(pad_gen3raw_input3),
	.pad_gen4raw_input(pad_gen4raw_input3),
	.pad_gen5raw_input(pad_gen5raw_input3),
	.pad_gen6raw_input(pad_gen6raw_input3),
	.pad_gen7raw_input(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out3),
	.phy_ddio_dmdout_0(phy_ddio_dmdout_0),
	.phy_ddio_dmdout_1(phy_ddio_dmdout_1),
	.phy_ddio_dmdout_2(phy_ddio_dmdout_2),
	.phy_ddio_dmdout_3(phy_ddio_dmdout_3),
	.phy_ddio_dqdout_0(phy_ddio_dqdout_0),
	.phy_ddio_dqdout_1(phy_ddio_dqdout_1),
	.phy_ddio_dqdout_2(phy_ddio_dqdout_2),
	.phy_ddio_dqdout_3(phy_ddio_dqdout_3),
	.phy_ddio_dqdout_4(phy_ddio_dqdout_4),
	.phy_ddio_dqdout_5(phy_ddio_dqdout_5),
	.phy_ddio_dqdout_6(phy_ddio_dqdout_6),
	.phy_ddio_dqdout_7(phy_ddio_dqdout_7),
	.phy_ddio_dqdout_8(phy_ddio_dqdout_8),
	.phy_ddio_dqdout_9(phy_ddio_dqdout_9),
	.phy_ddio_dqdout_10(phy_ddio_dqdout_10),
	.phy_ddio_dqdout_11(phy_ddio_dqdout_11),
	.phy_ddio_dqdout_12(phy_ddio_dqdout_12),
	.phy_ddio_dqdout_13(phy_ddio_dqdout_13),
	.phy_ddio_dqdout_14(phy_ddio_dqdout_14),
	.phy_ddio_dqdout_15(phy_ddio_dqdout_15),
	.phy_ddio_dqdout_16(phy_ddio_dqdout_16),
	.phy_ddio_dqdout_17(phy_ddio_dqdout_17),
	.phy_ddio_dqdout_18(phy_ddio_dqdout_18),
	.phy_ddio_dqdout_19(phy_ddio_dqdout_19),
	.phy_ddio_dqdout_20(phy_ddio_dqdout_20),
	.phy_ddio_dqdout_21(phy_ddio_dqdout_21),
	.phy_ddio_dqdout_22(phy_ddio_dqdout_22),
	.phy_ddio_dqdout_23(phy_ddio_dqdout_23),
	.phy_ddio_dqdout_24(phy_ddio_dqdout_24),
	.phy_ddio_dqdout_25(phy_ddio_dqdout_25),
	.phy_ddio_dqdout_26(phy_ddio_dqdout_26),
	.phy_ddio_dqdout_27(phy_ddio_dqdout_27),
	.phy_ddio_dqdout_28(phy_ddio_dqdout_28),
	.phy_ddio_dqdout_29(phy_ddio_dqdout_29),
	.phy_ddio_dqdout_30(phy_ddio_dqdout_30),
	.phy_ddio_dqdout_31(phy_ddio_dqdout_31),
	.phy_ddio_dqoe_0(phy_ddio_dqoe_0),
	.phy_ddio_dqoe_1(phy_ddio_dqoe_1),
	.phy_ddio_dqoe_2(phy_ddio_dqoe_2),
	.phy_ddio_dqoe_3(phy_ddio_dqoe_3),
	.phy_ddio_dqoe_4(phy_ddio_dqoe_4),
	.phy_ddio_dqoe_5(phy_ddio_dqoe_5),
	.phy_ddio_dqoe_6(phy_ddio_dqoe_6),
	.phy_ddio_dqoe_7(phy_ddio_dqoe_7),
	.phy_ddio_dqoe_8(phy_ddio_dqoe_8),
	.phy_ddio_dqoe_9(phy_ddio_dqoe_9),
	.phy_ddio_dqoe_10(phy_ddio_dqoe_10),
	.phy_ddio_dqoe_11(phy_ddio_dqoe_11),
	.phy_ddio_dqoe_12(phy_ddio_dqoe_12),
	.phy_ddio_dqoe_13(phy_ddio_dqoe_13),
	.phy_ddio_dqoe_14(phy_ddio_dqoe_14),
	.phy_ddio_dqoe_15(phy_ddio_dqoe_15),
	.phy_ddio_dqs_dout_0(phy_ddio_dqs_dout_0),
	.phy_ddio_dqs_dout_1(phy_ddio_dqs_dout_1),
	.phy_ddio_dqs_dout_2(phy_ddio_dqs_dout_2),
	.phy_ddio_dqs_dout_3(phy_ddio_dqs_dout_3),
	.phy_ddio_dqslogic_aclr_fifoctrl_0(phy_ddio_dqslogic_aclr_fifoctrl_0),
	.phy_ddio_dqslogic_aclr_pstamble_0(phy_ddio_dqslogic_aclr_pstamble_0),
	.phy_ddio_dqslogic_dqsena_0(phy_ddio_dqslogic_dqsena_0),
	.phy_ddio_dqslogic_dqsena_1(phy_ddio_dqslogic_dqsena_1),
	.phy_ddio_dqslogic_fiforeset_0(phy_ddio_dqslogic_fiforeset_0),
	.phy_ddio_dqslogic_incrdataen_0(phy_ddio_dqslogic_incrdataen_0),
	.phy_ddio_dqslogic_incrdataen_1(phy_ddio_dqslogic_incrdataen_1),
	.phy_ddio_dqslogic_incwrptr_0(phy_ddio_dqslogic_incwrptr_0),
	.phy_ddio_dqslogic_incwrptr_1(phy_ddio_dqslogic_incwrptr_1),
	.phy_ddio_dqslogic_oct_0(phy_ddio_dqslogic_oct_0),
	.phy_ddio_dqslogic_oct_1(phy_ddio_dqslogic_oct_1),
	.phy_ddio_dqslogic_readlatency_0(phy_ddio_dqslogic_readlatency_0),
	.phy_ddio_dqslogic_readlatency_1(phy_ddio_dqslogic_readlatency_1),
	.phy_ddio_dqslogic_readlatency_2(phy_ddio_dqslogic_readlatency_2),
	.phy_ddio_dqslogic_readlatency_3(phy_ddio_dqslogic_readlatency_3),
	.phy_ddio_dqslogic_readlatency_4(phy_ddio_dqslogic_readlatency_4),
	.phy_ddio_dqs_oe_0(phy_ddio_dqs_oe_0),
	.phy_ddio_dqs_oe_1(phy_ddio_dqs_oe_1),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_0),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_1),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_2),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_3),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_0),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_1),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_2),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_3),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_0),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_1),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_2),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_3),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_0),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_1),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_2),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_3),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_0),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_1),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_2),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_3),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_0),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_1),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_2),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_3),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_0),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_1),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_2),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_3),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_0),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_1),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_2),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_3),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[0]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

Computer_System_hps_sdram_p0_acv_hard_addr_cmd_pads uaddr_cmd_pads(
	.afi_clk(afi_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.phy_ddio_address_0(phy_ddio_address_0),
	.phy_ddio_address_1(phy_ddio_address_1),
	.phy_ddio_address_2(phy_ddio_address_2),
	.phy_ddio_address_3(phy_ddio_address_3),
	.phy_ddio_address_4(phy_ddio_address_4),
	.phy_ddio_address_5(phy_ddio_address_5),
	.phy_ddio_address_6(phy_ddio_address_6),
	.phy_ddio_address_7(phy_ddio_address_7),
	.phy_ddio_address_8(phy_ddio_address_8),
	.phy_ddio_address_9(phy_ddio_address_9),
	.phy_ddio_address_10(phy_ddio_address_10),
	.phy_ddio_address_11(phy_ddio_address_11),
	.phy_ddio_address_12(phy_ddio_address_12),
	.phy_ddio_address_13(phy_ddio_address_13),
	.phy_ddio_address_14(phy_ddio_address_14),
	.phy_ddio_address_15(phy_ddio_address_15),
	.phy_ddio_address_16(phy_ddio_address_16),
	.phy_ddio_address_17(phy_ddio_address_17),
	.phy_ddio_address_18(phy_ddio_address_18),
	.phy_ddio_address_19(phy_ddio_address_19),
	.phy_ddio_address_20(phy_ddio_address_20),
	.phy_ddio_address_21(phy_ddio_address_21),
	.phy_ddio_address_22(phy_ddio_address_22),
	.phy_ddio_address_23(phy_ddio_address_23),
	.phy_ddio_address_24(phy_ddio_address_24),
	.phy_ddio_address_25(phy_ddio_address_25),
	.phy_ddio_address_26(phy_ddio_address_26),
	.phy_ddio_address_27(phy_ddio_address_27),
	.phy_ddio_address_28(phy_ddio_address_28),
	.phy_ddio_address_29(phy_ddio_address_29),
	.phy_ddio_address_30(phy_ddio_address_30),
	.phy_ddio_address_31(phy_ddio_address_31),
	.phy_ddio_address_32(phy_ddio_address_32),
	.phy_ddio_address_33(phy_ddio_address_33),
	.phy_ddio_address_34(phy_ddio_address_34),
	.phy_ddio_address_35(phy_ddio_address_35),
	.phy_ddio_address_36(phy_ddio_address_36),
	.phy_ddio_address_37(phy_ddio_address_37),
	.phy_ddio_address_38(phy_ddio_address_38),
	.phy_ddio_address_39(phy_ddio_address_39),
	.phy_ddio_address_40(phy_ddio_address_40),
	.phy_ddio_address_41(phy_ddio_address_41),
	.phy_ddio_address_42(phy_ddio_address_42),
	.phy_ddio_address_43(phy_ddio_address_43),
	.phy_ddio_address_44(phy_ddio_address_44),
	.phy_ddio_address_45(phy_ddio_address_45),
	.phy_ddio_address_46(phy_ddio_address_46),
	.phy_ddio_address_47(phy_ddio_address_47),
	.phy_ddio_address_48(phy_ddio_address_48),
	.phy_ddio_address_49(phy_ddio_address_49),
	.phy_ddio_address_50(phy_ddio_address_50),
	.phy_ddio_address_51(phy_ddio_address_51),
	.phy_ddio_address_52(phy_ddio_address_52),
	.phy_ddio_address_53(phy_ddio_address_53),
	.phy_ddio_address_54(phy_ddio_address_54),
	.phy_ddio_address_55(phy_ddio_address_55),
	.phy_ddio_address_56(phy_ddio_address_56),
	.phy_ddio_address_57(phy_ddio_address_57),
	.phy_ddio_address_58(phy_ddio_address_58),
	.phy_ddio_address_59(phy_ddio_address_59),
	.phy_ddio_bank_0(phy_ddio_bank_0),
	.phy_ddio_bank_1(phy_ddio_bank_1),
	.phy_ddio_bank_2(phy_ddio_bank_2),
	.phy_ddio_bank_3(phy_ddio_bank_3),
	.phy_ddio_bank_4(phy_ddio_bank_4),
	.phy_ddio_bank_5(phy_ddio_bank_5),
	.phy_ddio_bank_6(phy_ddio_bank_6),
	.phy_ddio_bank_7(phy_ddio_bank_7),
	.phy_ddio_bank_8(phy_ddio_bank_8),
	.phy_ddio_bank_9(phy_ddio_bank_9),
	.phy_ddio_bank_10(phy_ddio_bank_10),
	.phy_ddio_bank_11(phy_ddio_bank_11),
	.phy_ddio_cas_n_0(phy_ddio_cas_n_0),
	.phy_ddio_cas_n_1(phy_ddio_cas_n_1),
	.phy_ddio_cas_n_2(phy_ddio_cas_n_2),
	.phy_ddio_cas_n_3(phy_ddio_cas_n_3),
	.phy_ddio_ck_0(phy_ddio_ck_0),
	.phy_ddio_ck_1(phy_ddio_ck_1),
	.phy_ddio_cke_0(phy_ddio_cke_0),
	.phy_ddio_cke_1(phy_ddio_cke_1),
	.phy_ddio_cke_2(phy_ddio_cke_2),
	.phy_ddio_cke_3(phy_ddio_cke_3),
	.phy_ddio_cs_n_0(phy_ddio_cs_n_0),
	.phy_ddio_cs_n_1(phy_ddio_cs_n_1),
	.phy_ddio_cs_n_2(phy_ddio_cs_n_2),
	.phy_ddio_cs_n_3(phy_ddio_cs_n_3),
	.phy_ddio_odt_0(phy_ddio_odt_0),
	.phy_ddio_odt_1(phy_ddio_odt_1),
	.phy_ddio_odt_2(phy_ddio_odt_2),
	.phy_ddio_odt_3(phy_ddio_odt_3),
	.phy_ddio_ras_n_0(phy_ddio_ras_n_0),
	.phy_ddio_ras_n_1(phy_ddio_ras_n_1),
	.phy_ddio_ras_n_2(phy_ddio_ras_n_2),
	.phy_ddio_ras_n_3(phy_ddio_ras_n_3),
	.phy_ddio_reset_n_0(phy_ddio_reset_n_0),
	.phy_ddio_reset_n_1(phy_ddio_reset_n_1),
	.phy_ddio_reset_n_2(phy_ddio_reset_n_2),
	.phy_ddio_reset_n_3(phy_ddio_reset_n_3),
	.phy_ddio_we_n_0(phy_ddio_we_n_0),
	.phy_ddio_we_n_1(phy_ddio_we_n_1),
	.phy_ddio_we_n_2(phy_ddio_we_n_2),
	.phy_ddio_we_n_3(phy_ddio_we_n_3),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6));

endmodule

module Computer_System_hps_sdram_p0_acv_hard_addr_cmd_pads (
	afi_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	phy_ddio_address_0,
	phy_ddio_address_1,
	phy_ddio_address_2,
	phy_ddio_address_3,
	phy_ddio_address_4,
	phy_ddio_address_5,
	phy_ddio_address_6,
	phy_ddio_address_7,
	phy_ddio_address_8,
	phy_ddio_address_9,
	phy_ddio_address_10,
	phy_ddio_address_11,
	phy_ddio_address_12,
	phy_ddio_address_13,
	phy_ddio_address_14,
	phy_ddio_address_15,
	phy_ddio_address_16,
	phy_ddio_address_17,
	phy_ddio_address_18,
	phy_ddio_address_19,
	phy_ddio_address_20,
	phy_ddio_address_21,
	phy_ddio_address_22,
	phy_ddio_address_23,
	phy_ddio_address_24,
	phy_ddio_address_25,
	phy_ddio_address_26,
	phy_ddio_address_27,
	phy_ddio_address_28,
	phy_ddio_address_29,
	phy_ddio_address_30,
	phy_ddio_address_31,
	phy_ddio_address_32,
	phy_ddio_address_33,
	phy_ddio_address_34,
	phy_ddio_address_35,
	phy_ddio_address_36,
	phy_ddio_address_37,
	phy_ddio_address_38,
	phy_ddio_address_39,
	phy_ddio_address_40,
	phy_ddio_address_41,
	phy_ddio_address_42,
	phy_ddio_address_43,
	phy_ddio_address_44,
	phy_ddio_address_45,
	phy_ddio_address_46,
	phy_ddio_address_47,
	phy_ddio_address_48,
	phy_ddio_address_49,
	phy_ddio_address_50,
	phy_ddio_address_51,
	phy_ddio_address_52,
	phy_ddio_address_53,
	phy_ddio_address_54,
	phy_ddio_address_55,
	phy_ddio_address_56,
	phy_ddio_address_57,
	phy_ddio_address_58,
	phy_ddio_address_59,
	phy_ddio_bank_0,
	phy_ddio_bank_1,
	phy_ddio_bank_2,
	phy_ddio_bank_3,
	phy_ddio_bank_4,
	phy_ddio_bank_5,
	phy_ddio_bank_6,
	phy_ddio_bank_7,
	phy_ddio_bank_8,
	phy_ddio_bank_9,
	phy_ddio_bank_10,
	phy_ddio_bank_11,
	phy_ddio_cas_n_0,
	phy_ddio_cas_n_1,
	phy_ddio_cas_n_2,
	phy_ddio_cas_n_3,
	phy_ddio_ck_0,
	phy_ddio_ck_1,
	phy_ddio_cke_0,
	phy_ddio_cke_1,
	phy_ddio_cke_2,
	phy_ddio_cke_3,
	phy_ddio_cs_n_0,
	phy_ddio_cs_n_1,
	phy_ddio_cs_n_2,
	phy_ddio_cs_n_3,
	phy_ddio_odt_0,
	phy_ddio_odt_1,
	phy_ddio_odt_2,
	phy_ddio_odt_3,
	phy_ddio_ras_n_0,
	phy_ddio_ras_n_1,
	phy_ddio_ras_n_2,
	phy_ddio_ras_n_3,
	phy_ddio_reset_n_0,
	phy_ddio_reset_n_1,
	phy_ddio_reset_n_2,
	phy_ddio_reset_n_3,
	phy_ddio_we_n_0,
	phy_ddio_we_n_1,
	phy_ddio_we_n_2,
	phy_ddio_we_n_3,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6)/* synthesis synthesis_greybox=0 */;
input 	afi_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	phy_ddio_address_0;
input 	phy_ddio_address_1;
input 	phy_ddio_address_2;
input 	phy_ddio_address_3;
input 	phy_ddio_address_4;
input 	phy_ddio_address_5;
input 	phy_ddio_address_6;
input 	phy_ddio_address_7;
input 	phy_ddio_address_8;
input 	phy_ddio_address_9;
input 	phy_ddio_address_10;
input 	phy_ddio_address_11;
input 	phy_ddio_address_12;
input 	phy_ddio_address_13;
input 	phy_ddio_address_14;
input 	phy_ddio_address_15;
input 	phy_ddio_address_16;
input 	phy_ddio_address_17;
input 	phy_ddio_address_18;
input 	phy_ddio_address_19;
input 	phy_ddio_address_20;
input 	phy_ddio_address_21;
input 	phy_ddio_address_22;
input 	phy_ddio_address_23;
input 	phy_ddio_address_24;
input 	phy_ddio_address_25;
input 	phy_ddio_address_26;
input 	phy_ddio_address_27;
input 	phy_ddio_address_28;
input 	phy_ddio_address_29;
input 	phy_ddio_address_30;
input 	phy_ddio_address_31;
input 	phy_ddio_address_32;
input 	phy_ddio_address_33;
input 	phy_ddio_address_34;
input 	phy_ddio_address_35;
input 	phy_ddio_address_36;
input 	phy_ddio_address_37;
input 	phy_ddio_address_38;
input 	phy_ddio_address_39;
input 	phy_ddio_address_40;
input 	phy_ddio_address_41;
input 	phy_ddio_address_42;
input 	phy_ddio_address_43;
input 	phy_ddio_address_44;
input 	phy_ddio_address_45;
input 	phy_ddio_address_46;
input 	phy_ddio_address_47;
input 	phy_ddio_address_48;
input 	phy_ddio_address_49;
input 	phy_ddio_address_50;
input 	phy_ddio_address_51;
input 	phy_ddio_address_52;
input 	phy_ddio_address_53;
input 	phy_ddio_address_54;
input 	phy_ddio_address_55;
input 	phy_ddio_address_56;
input 	phy_ddio_address_57;
input 	phy_ddio_address_58;
input 	phy_ddio_address_59;
input 	phy_ddio_bank_0;
input 	phy_ddio_bank_1;
input 	phy_ddio_bank_2;
input 	phy_ddio_bank_3;
input 	phy_ddio_bank_4;
input 	phy_ddio_bank_5;
input 	phy_ddio_bank_6;
input 	phy_ddio_bank_7;
input 	phy_ddio_bank_8;
input 	phy_ddio_bank_9;
input 	phy_ddio_bank_10;
input 	phy_ddio_bank_11;
input 	phy_ddio_cas_n_0;
input 	phy_ddio_cas_n_1;
input 	phy_ddio_cas_n_2;
input 	phy_ddio_cas_n_3;
input 	phy_ddio_ck_0;
input 	phy_ddio_ck_1;
input 	phy_ddio_cke_0;
input 	phy_ddio_cke_1;
input 	phy_ddio_cke_2;
input 	phy_ddio_cke_3;
input 	phy_ddio_cs_n_0;
input 	phy_ddio_cs_n_1;
input 	phy_ddio_cs_n_2;
input 	phy_ddio_cs_n_3;
input 	phy_ddio_odt_0;
input 	phy_ddio_odt_1;
input 	phy_ddio_odt_2;
input 	phy_ddio_odt_3;
input 	phy_ddio_ras_n_0;
input 	phy_ddio_ras_n_1;
input 	phy_ddio_ras_n_2;
input 	phy_ddio_ras_n_3;
input 	phy_ddio_reset_n_0;
input 	phy_ddio_reset_n_1;
input 	phy_ddio_reset_n_2;
input 	phy_ddio_reset_n_3;
input 	phy_ddio_we_n_0;
input 	phy_ddio_we_n_1;
input 	phy_ddio_we_n_2;
input 	phy_ddio_we_n_3;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \address_gen[0].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[1].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[2].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[3].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[4].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[5].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[6].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[7].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[8].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[9].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[10].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[11].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[12].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[13].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[14].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[15].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[16].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[17].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[19].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[18].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[21].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[22].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[23].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[24].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[20].acv_ac_ldc|adc_clk_cps ;
wire \clock_gen[0].umem_ck_pad|auto_generated|dataout[0] ;
wire \mem_ck_source[0] ;
wire \clock_gen[0].leveled_dqs_clocks[0] ;
wire \clock_gen[0].leveled_dqs_clocks[1] ;
wire \clock_gen[0].leveled_dqs_clocks[2] ;
wire \clock_gen[0].leveled_dqs_clocks[3] ;

wire [3:0] \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus ;

assign \clock_gen[0].leveled_dqs_clocks[0]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [0];
assign \clock_gen[0].leveled_dqs_clocks[1]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [1];
assign \clock_gen[0].leveled_dqs_clocks[2]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [2];
assign \clock_gen[0].leveled_dqs_clocks[3]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [3];

Computer_System_hps_sdram_p0_clock_pair_generator \clock_gen[0].uclk_generator (
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.datain({\clock_gen[0].umem_ck_pad|auto_generated|dataout[0] }));

Computer_System_altddio_out_1 \clock_gen[0].umem_ck_pad (
	.dataout({\clock_gen[0].umem_ck_pad|auto_generated|dataout[0] }),
	.datain_h({phy_ddio_ck_0}),
	.datain_l({phy_ddio_ck_1}),
	.outclock(\mem_ck_source[0] ));

Computer_System_hps_sdram_p0_generic_ddio_3 ureset_n_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk}),
	.dataout({dataout_unconnected_wire_14,dataout_unconnected_wire_13,dataout_unconnected_wire_12,dataout_unconnected_wire_11,dataout_unconnected_wire_10,dataout_unconnected_wire_9,dataout_unconnected_wire_8,dataout_unconnected_wire_7,dataout_unconnected_wire_6,
dataout_unconnected_wire_5,dataout_unconnected_wire_4,dataout_unconnected_wire_3,dataout_unconnected_wire_2,dataout_unconnected_wire_1,dataout_03}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[24].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_reset_n_3,phy_ddio_reset_n_2,phy_ddio_reset_n_1,phy_ddio_reset_n_0}));

Computer_System_hps_sdram_p0_generic_ddio_2 ucmd_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_unconnected_wire_14_1,dataout_unconnected_wire_13_1,dataout_unconnected_wire_12_1,dataout_unconnected_wire_11_1,dataout_unconnected_wire_10_1,dataout_unconnected_wire_9_1,dataout_unconnected_wire_8_1,dataout_unconnected_wire_7_1,
dataout_unconnected_wire_6_1,dataout_51,dataout_41,dataout_31,dataout_22,dataout_16,dataout_02}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[23].acv_ac_ldc|adc_clk_cps ,\address_gen[22].acv_ac_ldc|adc_clk_cps ,\address_gen[21].acv_ac_ldc|adc_clk_cps ,\address_gen[20].acv_ac_ldc|adc_clk_cps ,\address_gen[19].acv_ac_ldc|adc_clk_cps ,
\address_gen[18].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_we_n_3,phy_ddio_we_n_2,phy_ddio_we_n_1,phy_ddio_we_n_0,phy_ddio_cas_n_3,phy_ddio_cas_n_2,phy_ddio_cas_n_1,phy_ddio_cas_n_0,phy_ddio_ras_n_3,
phy_ddio_ras_n_2,phy_ddio_ras_n_1,phy_ddio_ras_n_0,phy_ddio_odt_3,phy_ddio_odt_2,phy_ddio_odt_1,phy_ddio_odt_0,phy_ddio_cke_3,phy_ddio_cke_2,phy_ddio_cke_1,phy_ddio_cke_0,phy_ddio_cs_n_3,phy_ddio_cs_n_2,phy_ddio_cs_n_1,phy_ddio_cs_n_0}));

Computer_System_hps_sdram_p0_generic_ddio_1 ubank_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_unconnected_wire_14_2,dataout_unconnected_wire_13_2,dataout_unconnected_wire_12_2,dataout_unconnected_wire_11_2,dataout_unconnected_wire_10_2,dataout_unconnected_wire_9_2,dataout_unconnected_wire_8_2,dataout_unconnected_wire_7_2,
dataout_unconnected_wire_6_2,dataout_unconnected_wire_5_1,dataout_unconnected_wire_4_1,dataout_unconnected_wire_3_1,dataout_21,dataout_15,dataout_01}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[17].acv_ac_ldc|adc_clk_cps ,\address_gen[16].acv_ac_ldc|adc_clk_cps ,\address_gen[15].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_bank_11,phy_ddio_bank_10,phy_ddio_bank_9,phy_ddio_bank_8,phy_ddio_bank_7,phy_ddio_bank_6,phy_ddio_bank_5,
phy_ddio_bank_4,phy_ddio_bank_3,phy_ddio_bank_2,phy_ddio_bank_1,phy_ddio_bank_0}));

Computer_System_hps_sdram_p0_generic_ddio uaddress_pad(
	.clk_hr({afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_14,dataout_13,dataout_12,dataout_11,dataout_10,dataout_9,dataout_8,dataout_7,dataout_6,dataout_5,dataout_4,dataout_3,dataout_2,dataout_1,dataout_0}),
	.clk_fr({\address_gen[14].acv_ac_ldc|adc_clk_cps ,\address_gen[13].acv_ac_ldc|adc_clk_cps ,\address_gen[12].acv_ac_ldc|adc_clk_cps ,\address_gen[11].acv_ac_ldc|adc_clk_cps ,\address_gen[10].acv_ac_ldc|adc_clk_cps ,\address_gen[9].acv_ac_ldc|adc_clk_cps ,
\address_gen[8].acv_ac_ldc|adc_clk_cps ,\address_gen[7].acv_ac_ldc|adc_clk_cps ,\address_gen[6].acv_ac_ldc|adc_clk_cps ,\address_gen[5].acv_ac_ldc|adc_clk_cps ,\address_gen[4].acv_ac_ldc|adc_clk_cps ,\address_gen[3].acv_ac_ldc|adc_clk_cps ,
\address_gen[2].acv_ac_ldc|adc_clk_cps ,\address_gen[1].acv_ac_ldc|adc_clk_cps ,\address_gen[0].acv_ac_ldc|adc_clk_cps }),
	.datain({phy_ddio_address_59,phy_ddio_address_58,phy_ddio_address_57,phy_ddio_address_56,phy_ddio_address_55,phy_ddio_address_54,phy_ddio_address_53,phy_ddio_address_52,phy_ddio_address_51,phy_ddio_address_50,phy_ddio_address_49,phy_ddio_address_48,phy_ddio_address_47,
phy_ddio_address_46,phy_ddio_address_45,phy_ddio_address_44,phy_ddio_address_43,phy_ddio_address_42,phy_ddio_address_41,phy_ddio_address_40,phy_ddio_address_39,phy_ddio_address_38,phy_ddio_address_37,phy_ddio_address_36,phy_ddio_address_35,phy_ddio_address_34,
phy_ddio_address_33,phy_ddio_address_32,phy_ddio_address_31,phy_ddio_address_30,phy_ddio_address_29,phy_ddio_address_28,phy_ddio_address_27,phy_ddio_address_26,phy_ddio_address_25,phy_ddio_address_24,phy_ddio_address_23,phy_ddio_address_22,phy_ddio_address_21,
phy_ddio_address_20,phy_ddio_address_19,phy_ddio_address_18,phy_ddio_address_17,phy_ddio_address_16,phy_ddio_address_15,phy_ddio_address_14,phy_ddio_address_13,phy_ddio_address_12,phy_ddio_address_11,phy_ddio_address_10,phy_ddio_address_9,phy_ddio_address_8,
phy_ddio_address_7,phy_ddio_address_6,phy_ddio_address_5,phy_ddio_address_4,phy_ddio_address_3,phy_ddio_address_2,phy_ddio_address_1,phy_ddio_address_0}));

Computer_System_hps_sdram_p0_acv_ldc_16 \address_gen[24].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[24].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_15 \address_gen[23].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[23].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_14 \address_gen[22].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[22].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_13 \address_gen[21].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[21].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_12 \address_gen[20].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[20].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_10 \address_gen[19].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[19].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_9 \address_gen[18].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[18].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_8 \address_gen[17].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[17].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_7 \address_gen[16].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[16].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_6 \address_gen[15].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[15].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_5 \address_gen[14].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[14].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_4 \address_gen[13].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[13].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_3 \address_gen[12].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[12].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_2 \address_gen[11].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[11].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_1 \address_gen[10].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[10].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_24 \address_gen[9].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[9].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_23 \address_gen[8].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[8].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_22 \address_gen[7].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[7].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_21 \address_gen[6].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[6].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_20 \address_gen[5].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[5].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_19 \address_gen[4].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[4].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_18 \address_gen[3].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[3].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_17 \address_gen[2].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[2].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc_11 \address_gen[1].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[1].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

Computer_System_hps_sdram_p0_acv_ldc \address_gen[0].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[0].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

cyclonev_clk_phase_select \clock_gen[0].clk_phase_select_dqs (
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\clock_gen[0].leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(\mem_ck_source[0] ));
defparam \clock_gen[0].clk_phase_select_dqs .invert_phase = "false";
defparam \clock_gen[0].clk_phase_select_dqs .phase_setting = 0;
defparam \clock_gen[0].clk_phase_select_dqs .physical_clock_source = "dqs";
defparam \clock_gen[0].clk_phase_select_dqs .use_dqs_input = "false";
defparam \clock_gen[0].clk_phase_select_dqs .use_phasectrlin = "false";

cyclonev_leveling_delay_chain \clock_gen[0].leveling_delay_chain_dqs (
	.clkin(afi_clk),
	.delayctrlin({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.clkout(\clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus ));
defparam \clock_gen[0].leveling_delay_chain_dqs .physical_clock_source = "dqs";
defparam \clock_gen[0].leveling_delay_chain_dqs .sim_buffer_delay_increment = 10;
defparam \clock_gen[0].leveling_delay_chain_dqs .sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_altddio_out_1 (
	dataout,
	datain_h,
	datain_l,
	outclock)/* synthesis synthesis_greybox=0 */;
inout 	[0:0] dataout;
input 	[0:0] datain_h;
input 	[0:0] datain_l;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_ddio_out_uqe auto_generated(
	.dataout({dataout[0]}),
	.datain_h({datain_h[0]}),
	.datain_l({datain_l[0]}),
	.outclock(outclock));

endmodule

module Computer_System_ddio_out_uqe (
	dataout,
	datain_h,
	datain_l,
	outclock)/* synthesis synthesis_greybox=0 */;
output 	[0:0] dataout;
input 	[0:0] datain_h;
input 	[0:0] datain_l;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "none";
defparam \ddio_outa[0] .half_rate_mode = "false";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_acv_ldc (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_1 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_2 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_3 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_4 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_5 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_6 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_7 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_8 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_9 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_10 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_11 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_12 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_13 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_14 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_15 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_16 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_17 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_18 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_19 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_20 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_21 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_22 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_23 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_24 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_p0_clock_pair_generator (
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	datain)/* synthesis synthesis_greybox=0 */;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	[0:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(datain[0]),
	.oein(gnd),
	.dtcin(gnd),
	.o(wire_pseudo_diffa_o_0),
	.obar(wire_pseudo_diffa_obar_0),
	.oeout(wire_pseudo_diffa_oeout_0),
	.oebout(wire_pseudo_diffa_oebout_0),
	.dtc(),
	.dtcbar());

endmodule

module Computer_System_hps_sdram_p0_generic_ddio (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;
wire \acblock[3].fr_data_lo ;
wire \acblock[3].fr_data_hi ;
wire \acblock[4].fr_data_lo ;
wire \acblock[4].fr_data_hi ;
wire \acblock[5].fr_data_lo ;
wire \acblock[5].fr_data_hi ;
wire \acblock[6].fr_data_lo ;
wire \acblock[6].fr_data_hi ;
wire \acblock[7].fr_data_lo ;
wire \acblock[7].fr_data_hi ;
wire \acblock[8].fr_data_lo ;
wire \acblock[8].fr_data_hi ;
wire \acblock[9].fr_data_lo ;
wire \acblock[9].fr_data_hi ;
wire \acblock[10].fr_data_lo ;
wire \acblock[10].fr_data_hi ;
wire \acblock[11].fr_data_lo ;
wire \acblock[11].fr_data_hi ;
wire \acblock[12].fr_data_lo ;
wire \acblock[12].fr_data_hi ;
wire \acblock[13].fr_data_lo ;
wire \acblock[13].fr_data_hi ;
wire \acblock[14].fr_data_lo ;
wire \acblock[14].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].ddio_out (
	.datainlo(\acblock[3].fr_data_lo ),
	.datainhi(\acblock[3].fr_data_hi ),
	.clkhi(clk_fr[3]),
	.clklo(clk_fr[3]),
	.muxsel(clk_fr[3]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[3]),
	.dfflo(),
	.dffhi());
defparam \acblock[3].ddio_out .async_mode = "none";
defparam \acblock[3].ddio_out .half_rate_mode = "false";
defparam \acblock[3].ddio_out .power_up = "low";
defparam \acblock[3].ddio_out .sync_mode = "none";
defparam \acblock[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].ddio_out (
	.datainlo(\acblock[4].fr_data_lo ),
	.datainhi(\acblock[4].fr_data_hi ),
	.clkhi(clk_fr[4]),
	.clklo(clk_fr[4]),
	.muxsel(clk_fr[4]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[4]),
	.dfflo(),
	.dffhi());
defparam \acblock[4].ddio_out .async_mode = "none";
defparam \acblock[4].ddio_out .half_rate_mode = "false";
defparam \acblock[4].ddio_out .power_up = "low";
defparam \acblock[4].ddio_out .sync_mode = "none";
defparam \acblock[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].ddio_out (
	.datainlo(\acblock[5].fr_data_lo ),
	.datainhi(\acblock[5].fr_data_hi ),
	.clkhi(clk_fr[5]),
	.clklo(clk_fr[5]),
	.muxsel(clk_fr[5]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[5]),
	.dfflo(),
	.dffhi());
defparam \acblock[5].ddio_out .async_mode = "none";
defparam \acblock[5].ddio_out .half_rate_mode = "false";
defparam \acblock[5].ddio_out .power_up = "low";
defparam \acblock[5].ddio_out .sync_mode = "none";
defparam \acblock[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].ddio_out (
	.datainlo(\acblock[6].fr_data_lo ),
	.datainhi(\acblock[6].fr_data_hi ),
	.clkhi(clk_fr[6]),
	.clklo(clk_fr[6]),
	.muxsel(clk_fr[6]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[6]),
	.dfflo(),
	.dffhi());
defparam \acblock[6].ddio_out .async_mode = "none";
defparam \acblock[6].ddio_out .half_rate_mode = "false";
defparam \acblock[6].ddio_out .power_up = "low";
defparam \acblock[6].ddio_out .sync_mode = "none";
defparam \acblock[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].ddio_out (
	.datainlo(\acblock[7].fr_data_lo ),
	.datainhi(\acblock[7].fr_data_hi ),
	.clkhi(clk_fr[7]),
	.clklo(clk_fr[7]),
	.muxsel(clk_fr[7]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[7]),
	.dfflo(),
	.dffhi());
defparam \acblock[7].ddio_out .async_mode = "none";
defparam \acblock[7].ddio_out .half_rate_mode = "false";
defparam \acblock[7].ddio_out .power_up = "low";
defparam \acblock[7].ddio_out .sync_mode = "none";
defparam \acblock[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].ddio_out (
	.datainlo(\acblock[8].fr_data_lo ),
	.datainhi(\acblock[8].fr_data_hi ),
	.clkhi(clk_fr[8]),
	.clklo(clk_fr[8]),
	.muxsel(clk_fr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[8]),
	.dfflo(),
	.dffhi());
defparam \acblock[8].ddio_out .async_mode = "none";
defparam \acblock[8].ddio_out .half_rate_mode = "false";
defparam \acblock[8].ddio_out .power_up = "low";
defparam \acblock[8].ddio_out .sync_mode = "none";
defparam \acblock[8].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].ddio_out (
	.datainlo(\acblock[9].fr_data_lo ),
	.datainhi(\acblock[9].fr_data_hi ),
	.clkhi(clk_fr[9]),
	.clklo(clk_fr[9]),
	.muxsel(clk_fr[9]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[9]),
	.dfflo(),
	.dffhi());
defparam \acblock[9].ddio_out .async_mode = "none";
defparam \acblock[9].ddio_out .half_rate_mode = "false";
defparam \acblock[9].ddio_out .power_up = "low";
defparam \acblock[9].ddio_out .sync_mode = "none";
defparam \acblock[9].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].ddio_out (
	.datainlo(\acblock[10].fr_data_lo ),
	.datainhi(\acblock[10].fr_data_hi ),
	.clkhi(clk_fr[10]),
	.clklo(clk_fr[10]),
	.muxsel(clk_fr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[10]),
	.dfflo(),
	.dffhi());
defparam \acblock[10].ddio_out .async_mode = "none";
defparam \acblock[10].ddio_out .half_rate_mode = "false";
defparam \acblock[10].ddio_out .power_up = "low";
defparam \acblock[10].ddio_out .sync_mode = "none";
defparam \acblock[10].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].ddio_out (
	.datainlo(\acblock[11].fr_data_lo ),
	.datainhi(\acblock[11].fr_data_hi ),
	.clkhi(clk_fr[11]),
	.clklo(clk_fr[11]),
	.muxsel(clk_fr[11]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[11]),
	.dfflo(),
	.dffhi());
defparam \acblock[11].ddio_out .async_mode = "none";
defparam \acblock[11].ddio_out .half_rate_mode = "false";
defparam \acblock[11].ddio_out .power_up = "low";
defparam \acblock[11].ddio_out .sync_mode = "none";
defparam \acblock[11].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].ddio_out (
	.datainlo(\acblock[12].fr_data_lo ),
	.datainhi(\acblock[12].fr_data_hi ),
	.clkhi(clk_fr[12]),
	.clklo(clk_fr[12]),
	.muxsel(clk_fr[12]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[12]),
	.dfflo(),
	.dffhi());
defparam \acblock[12].ddio_out .async_mode = "none";
defparam \acblock[12].ddio_out .half_rate_mode = "false";
defparam \acblock[12].ddio_out .power_up = "low";
defparam \acblock[12].ddio_out .sync_mode = "none";
defparam \acblock[12].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].ddio_out (
	.datainlo(\acblock[13].fr_data_lo ),
	.datainhi(\acblock[13].fr_data_hi ),
	.clkhi(clk_fr[13]),
	.clklo(clk_fr[13]),
	.muxsel(clk_fr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[13]),
	.dfflo(),
	.dffhi());
defparam \acblock[13].ddio_out .async_mode = "none";
defparam \acblock[13].ddio_out .half_rate_mode = "false";
defparam \acblock[13].ddio_out .power_up = "low";
defparam \acblock[13].ddio_out .sync_mode = "none";
defparam \acblock[13].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].ddio_out (
	.datainlo(\acblock[14].fr_data_lo ),
	.datainhi(\acblock[14].fr_data_hi ),
	.clkhi(clk_fr[14]),
	.clklo(clk_fr[14]),
	.muxsel(clk_fr[14]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[14]),
	.dfflo(),
	.dffhi());
defparam \acblock[14].ddio_out .async_mode = "none";
defparam \acblock[14].ddio_out .half_rate_mode = "false";
defparam \acblock[14].ddio_out .power_up = "low";
defparam \acblock[14].ddio_out .sync_mode = "none";
defparam \acblock[14].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_lo (
	.datainlo(datain[15]),
	.datainhi(datain[13]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_lo .async_mode = "none";
defparam \acblock[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_lo .power_up = "low";
defparam \acblock[3].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_hi (
	.datainlo(datain[14]),
	.datainhi(datain[12]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_hi .async_mode = "none";
defparam \acblock[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_hi .power_up = "low";
defparam \acblock[3].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_lo (
	.datainlo(datain[19]),
	.datainhi(datain[17]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_lo .async_mode = "none";
defparam \acblock[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_lo .power_up = "low";
defparam \acblock[4].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_hi (
	.datainlo(datain[18]),
	.datainhi(datain[16]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_hi .async_mode = "none";
defparam \acblock[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_hi .power_up = "low";
defparam \acblock[4].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_lo (
	.datainlo(datain[23]),
	.datainhi(datain[21]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_lo .async_mode = "none";
defparam \acblock[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_lo .power_up = "low";
defparam \acblock[5].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_hi (
	.datainlo(datain[22]),
	.datainhi(datain[20]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_hi .async_mode = "none";
defparam \acblock[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_hi .power_up = "low";
defparam \acblock[5].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].hr_to_fr_lo (
	.datainlo(datain[27]),
	.datainhi(datain[25]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[6].hr_to_fr_lo .async_mode = "none";
defparam \acblock[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[6].hr_to_fr_lo .power_up = "low";
defparam \acblock[6].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].hr_to_fr_hi (
	.datainlo(datain[26]),
	.datainhi(datain[24]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[6].hr_to_fr_hi .async_mode = "none";
defparam \acblock[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[6].hr_to_fr_hi .power_up = "low";
defparam \acblock[6].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].hr_to_fr_lo (
	.datainlo(datain[31]),
	.datainhi(datain[29]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[7].hr_to_fr_lo .async_mode = "none";
defparam \acblock[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[7].hr_to_fr_lo .power_up = "low";
defparam \acblock[7].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].hr_to_fr_hi (
	.datainlo(datain[30]),
	.datainhi(datain[28]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[7].hr_to_fr_hi .async_mode = "none";
defparam \acblock[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[7].hr_to_fr_hi .power_up = "low";
defparam \acblock[7].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].hr_to_fr_lo (
	.datainlo(datain[35]),
	.datainhi(datain[33]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[8].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[8].hr_to_fr_lo .async_mode = "none";
defparam \acblock[8].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[8].hr_to_fr_lo .power_up = "low";
defparam \acblock[8].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[8].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].hr_to_fr_hi (
	.datainlo(datain[34]),
	.datainhi(datain[32]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[8].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[8].hr_to_fr_hi .async_mode = "none";
defparam \acblock[8].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[8].hr_to_fr_hi .power_up = "low";
defparam \acblock[8].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[8].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].hr_to_fr_lo (
	.datainlo(datain[39]),
	.datainhi(datain[37]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[9].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[9].hr_to_fr_lo .async_mode = "none";
defparam \acblock[9].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[9].hr_to_fr_lo .power_up = "low";
defparam \acblock[9].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[9].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].hr_to_fr_hi (
	.datainlo(datain[38]),
	.datainhi(datain[36]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[9].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[9].hr_to_fr_hi .async_mode = "none";
defparam \acblock[9].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[9].hr_to_fr_hi .power_up = "low";
defparam \acblock[9].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[9].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].hr_to_fr_lo (
	.datainlo(datain[43]),
	.datainhi(datain[41]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[10].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[10].hr_to_fr_lo .async_mode = "none";
defparam \acblock[10].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[10].hr_to_fr_lo .power_up = "low";
defparam \acblock[10].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[10].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].hr_to_fr_hi (
	.datainlo(datain[42]),
	.datainhi(datain[40]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[10].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[10].hr_to_fr_hi .async_mode = "none";
defparam \acblock[10].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[10].hr_to_fr_hi .power_up = "low";
defparam \acblock[10].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[10].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].hr_to_fr_lo (
	.datainlo(datain[47]),
	.datainhi(datain[45]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[11].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[11].hr_to_fr_lo .async_mode = "none";
defparam \acblock[11].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[11].hr_to_fr_lo .power_up = "low";
defparam \acblock[11].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[11].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].hr_to_fr_hi (
	.datainlo(datain[46]),
	.datainhi(datain[44]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[11].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[11].hr_to_fr_hi .async_mode = "none";
defparam \acblock[11].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[11].hr_to_fr_hi .power_up = "low";
defparam \acblock[11].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[11].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].hr_to_fr_lo (
	.datainlo(datain[51]),
	.datainhi(datain[49]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[12].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[12].hr_to_fr_lo .async_mode = "none";
defparam \acblock[12].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[12].hr_to_fr_lo .power_up = "low";
defparam \acblock[12].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[12].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].hr_to_fr_hi (
	.datainlo(datain[50]),
	.datainhi(datain[48]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[12].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[12].hr_to_fr_hi .async_mode = "none";
defparam \acblock[12].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[12].hr_to_fr_hi .power_up = "low";
defparam \acblock[12].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[12].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].hr_to_fr_lo (
	.datainlo(datain[55]),
	.datainhi(datain[53]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[13].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[13].hr_to_fr_lo .async_mode = "none";
defparam \acblock[13].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[13].hr_to_fr_lo .power_up = "low";
defparam \acblock[13].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[13].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].hr_to_fr_hi (
	.datainlo(datain[54]),
	.datainhi(datain[52]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[13].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[13].hr_to_fr_hi .async_mode = "none";
defparam \acblock[13].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[13].hr_to_fr_hi .power_up = "low";
defparam \acblock[13].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[13].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].hr_to_fr_lo (
	.datainlo(datain[59]),
	.datainhi(datain[57]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[14].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[14].hr_to_fr_lo .async_mode = "none";
defparam \acblock[14].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[14].hr_to_fr_lo .power_up = "low";
defparam \acblock[14].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[14].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].hr_to_fr_hi (
	.datainlo(datain[58]),
	.datainhi(datain[56]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[14].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[14].hr_to_fr_hi .async_mode = "none";
defparam \acblock[14].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[14].hr_to_fr_hi .power_up = "low";
defparam \acblock[14].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[14].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_generic_ddio_1 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_generic_ddio_2 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[3].fr_data_lo ;
wire \acblock[3].fr_data_hi ;
wire \acblock[4].fr_data_lo ;
wire \acblock[4].fr_data_hi ;
wire \acblock[5].fr_data_lo ;
wire \acblock[5].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;


cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].ddio_out (
	.datainlo(\acblock[3].fr_data_lo ),
	.datainhi(\acblock[3].fr_data_hi ),
	.clkhi(clk_fr[3]),
	.clklo(clk_fr[3]),
	.muxsel(clk_fr[3]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[3]),
	.dfflo(),
	.dffhi());
defparam \acblock[3].ddio_out .async_mode = "none";
defparam \acblock[3].ddio_out .half_rate_mode = "false";
defparam \acblock[3].ddio_out .power_up = "low";
defparam \acblock[3].ddio_out .sync_mode = "none";
defparam \acblock[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].ddio_out (
	.datainlo(\acblock[4].fr_data_lo ),
	.datainhi(\acblock[4].fr_data_hi ),
	.clkhi(clk_fr[4]),
	.clklo(clk_fr[4]),
	.muxsel(clk_fr[4]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[4]),
	.dfflo(),
	.dffhi());
defparam \acblock[4].ddio_out .async_mode = "none";
defparam \acblock[4].ddio_out .half_rate_mode = "false";
defparam \acblock[4].ddio_out .power_up = "low";
defparam \acblock[4].ddio_out .sync_mode = "none";
defparam \acblock[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].ddio_out (
	.datainlo(\acblock[5].fr_data_lo ),
	.datainhi(\acblock[5].fr_data_hi ),
	.clkhi(clk_fr[5]),
	.clklo(clk_fr[5]),
	.muxsel(clk_fr[5]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[5]),
	.dfflo(),
	.dffhi());
defparam \acblock[5].ddio_out .async_mode = "none";
defparam \acblock[5].ddio_out .half_rate_mode = "false";
defparam \acblock[5].ddio_out .power_up = "low";
defparam \acblock[5].ddio_out .sync_mode = "none";
defparam \acblock[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_lo (
	.datainlo(datain[15]),
	.datainhi(datain[13]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_lo .async_mode = "none";
defparam \acblock[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_lo .power_up = "low";
defparam \acblock[3].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_hi (
	.datainlo(datain[14]),
	.datainhi(datain[12]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_hi .async_mode = "none";
defparam \acblock[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_hi .power_up = "low";
defparam \acblock[3].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_lo (
	.datainlo(datain[19]),
	.datainhi(datain[17]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_lo .async_mode = "none";
defparam \acblock[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_lo .power_up = "low";
defparam \acblock[4].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_hi (
	.datainlo(datain[18]),
	.datainhi(datain[16]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_hi .async_mode = "none";
defparam \acblock[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_hi .power_up = "low";
defparam \acblock[4].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_lo (
	.datainlo(datain[23]),
	.datainhi(datain[21]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_lo .async_mode = "none";
defparam \acblock[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_lo .power_up = "low";
defparam \acblock[5].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_hi (
	.datainlo(datain[22]),
	.datainhi(datain[20]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_hi .async_mode = "none";
defparam \acblock[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_hi .power_up = "low";
defparam \acblock[5].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_generic_ddio_3 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_altdqdqs (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_0,
	phy_ddio_dmdout_1,
	phy_ddio_dmdout_2,
	phy_ddio_dmdout_3,
	phy_ddio_dqdout_0,
	phy_ddio_dqdout_1,
	phy_ddio_dqdout_2,
	phy_ddio_dqdout_3,
	phy_ddio_dqdout_4,
	phy_ddio_dqdout_5,
	phy_ddio_dqdout_6,
	phy_ddio_dqdout_7,
	phy_ddio_dqdout_8,
	phy_ddio_dqdout_9,
	phy_ddio_dqdout_10,
	phy_ddio_dqdout_11,
	phy_ddio_dqdout_12,
	phy_ddio_dqdout_13,
	phy_ddio_dqdout_14,
	phy_ddio_dqdout_15,
	phy_ddio_dqdout_16,
	phy_ddio_dqdout_17,
	phy_ddio_dqdout_18,
	phy_ddio_dqdout_19,
	phy_ddio_dqdout_20,
	phy_ddio_dqdout_21,
	phy_ddio_dqdout_22,
	phy_ddio_dqdout_23,
	phy_ddio_dqdout_24,
	phy_ddio_dqdout_25,
	phy_ddio_dqdout_26,
	phy_ddio_dqdout_27,
	phy_ddio_dqdout_28,
	phy_ddio_dqdout_29,
	phy_ddio_dqdout_30,
	phy_ddio_dqdout_31,
	phy_ddio_dqoe_0,
	phy_ddio_dqoe_1,
	phy_ddio_dqoe_2,
	phy_ddio_dqoe_3,
	phy_ddio_dqoe_4,
	phy_ddio_dqoe_5,
	phy_ddio_dqoe_6,
	phy_ddio_dqoe_7,
	phy_ddio_dqoe_8,
	phy_ddio_dqoe_9,
	phy_ddio_dqoe_10,
	phy_ddio_dqoe_11,
	phy_ddio_dqoe_12,
	phy_ddio_dqoe_13,
	phy_ddio_dqoe_14,
	phy_ddio_dqoe_15,
	phy_ddio_dqs_dout_0,
	phy_ddio_dqs_dout_1,
	phy_ddio_dqs_dout_2,
	phy_ddio_dqs_dout_3,
	phy_ddio_dqslogic_aclr_fifoctrl_0,
	phy_ddio_dqslogic_aclr_pstamble_0,
	phy_ddio_dqslogic_dqsena_0,
	phy_ddio_dqslogic_dqsena_1,
	phy_ddio_dqslogic_fiforeset_0,
	phy_ddio_dqslogic_incrdataen_0,
	phy_ddio_dqslogic_incrdataen_1,
	phy_ddio_dqslogic_incwrptr_0,
	phy_ddio_dqslogic_incwrptr_1,
	phy_ddio_dqslogic_oct_0,
	phy_ddio_dqslogic_oct_1,
	phy_ddio_dqslogic_readlatency_0,
	phy_ddio_dqslogic_readlatency_1,
	phy_ddio_dqslogic_readlatency_2,
	phy_ddio_dqslogic_readlatency_3,
	phy_ddio_dqslogic_readlatency_4,
	phy_ddio_dqs_oe_0,
	phy_ddio_dqs_oe_1,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_0;
input 	phy_ddio_dmdout_1;
input 	phy_ddio_dmdout_2;
input 	phy_ddio_dmdout_3;
input 	phy_ddio_dqdout_0;
input 	phy_ddio_dqdout_1;
input 	phy_ddio_dqdout_2;
input 	phy_ddio_dqdout_3;
input 	phy_ddio_dqdout_4;
input 	phy_ddio_dqdout_5;
input 	phy_ddio_dqdout_6;
input 	phy_ddio_dqdout_7;
input 	phy_ddio_dqdout_8;
input 	phy_ddio_dqdout_9;
input 	phy_ddio_dqdout_10;
input 	phy_ddio_dqdout_11;
input 	phy_ddio_dqdout_12;
input 	phy_ddio_dqdout_13;
input 	phy_ddio_dqdout_14;
input 	phy_ddio_dqdout_15;
input 	phy_ddio_dqdout_16;
input 	phy_ddio_dqdout_17;
input 	phy_ddio_dqdout_18;
input 	phy_ddio_dqdout_19;
input 	phy_ddio_dqdout_20;
input 	phy_ddio_dqdout_21;
input 	phy_ddio_dqdout_22;
input 	phy_ddio_dqdout_23;
input 	phy_ddio_dqdout_24;
input 	phy_ddio_dqdout_25;
input 	phy_ddio_dqdout_26;
input 	phy_ddio_dqdout_27;
input 	phy_ddio_dqdout_28;
input 	phy_ddio_dqdout_29;
input 	phy_ddio_dqdout_30;
input 	phy_ddio_dqdout_31;
input 	phy_ddio_dqoe_0;
input 	phy_ddio_dqoe_1;
input 	phy_ddio_dqoe_2;
input 	phy_ddio_dqoe_3;
input 	phy_ddio_dqoe_4;
input 	phy_ddio_dqoe_5;
input 	phy_ddio_dqoe_6;
input 	phy_ddio_dqoe_7;
input 	phy_ddio_dqoe_8;
input 	phy_ddio_dqoe_9;
input 	phy_ddio_dqoe_10;
input 	phy_ddio_dqoe_11;
input 	phy_ddio_dqoe_12;
input 	phy_ddio_dqoe_13;
input 	phy_ddio_dqoe_14;
input 	phy_ddio_dqoe_15;
input 	phy_ddio_dqs_dout_0;
input 	phy_ddio_dqs_dout_1;
input 	phy_ddio_dqs_dout_2;
input 	phy_ddio_dqs_dout_3;
input 	phy_ddio_dqslogic_aclr_fifoctrl_0;
input 	phy_ddio_dqslogic_aclr_pstamble_0;
input 	phy_ddio_dqslogic_dqsena_0;
input 	phy_ddio_dqslogic_dqsena_1;
input 	phy_ddio_dqslogic_fiforeset_0;
input 	phy_ddio_dqslogic_incrdataen_0;
input 	phy_ddio_dqslogic_incrdataen_1;
input 	phy_ddio_dqslogic_incwrptr_0;
input 	phy_ddio_dqslogic_incwrptr_1;
input 	phy_ddio_dqslogic_oct_0;
input 	phy_ddio_dqslogic_oct_1;
input 	phy_ddio_dqslogic_readlatency_0;
input 	phy_ddio_dqslogic_readlatency_1;
input 	phy_ddio_dqslogic_readlatency_2;
input 	phy_ddio_dqslogic_readlatency_3;
input 	phy_ddio_dqslogic_readlatency_4;
input 	phy_ddio_dqs_oe_0;
input 	phy_ddio_dqs_oe_1;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.config_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_3,phy_ddio_dmdout_2,phy_ddio_dmdout_1,phy_ddio_dmdout_0}),
	.write_data_in({phy_ddio_dqdout_31,phy_ddio_dqdout_30,phy_ddio_dqdout_29,phy_ddio_dqdout_28,phy_ddio_dqdout_27,phy_ddio_dqdout_26,phy_ddio_dqdout_25,phy_ddio_dqdout_24,phy_ddio_dqdout_23,phy_ddio_dqdout_22,phy_ddio_dqdout_21,phy_ddio_dqdout_20,phy_ddio_dqdout_19,phy_ddio_dqdout_18,
phy_ddio_dqdout_17,phy_ddio_dqdout_16,phy_ddio_dqdout_15,phy_ddio_dqdout_14,phy_ddio_dqdout_13,phy_ddio_dqdout_12,phy_ddio_dqdout_11,phy_ddio_dqdout_10,phy_ddio_dqdout_9,phy_ddio_dqdout_8,phy_ddio_dqdout_7,phy_ddio_dqdout_6,phy_ddio_dqdout_5,phy_ddio_dqdout_4,
phy_ddio_dqdout_3,phy_ddio_dqdout_2,phy_ddio_dqdout_1,phy_ddio_dqdout_0}),
	.write_oe_in({phy_ddio_dqoe_15,phy_ddio_dqoe_14,phy_ddio_dqoe_13,phy_ddio_dqoe_12,phy_ddio_dqoe_11,phy_ddio_dqoe_10,phy_ddio_dqoe_9,phy_ddio_dqoe_8,phy_ddio_dqoe_7,phy_ddio_dqoe_6,phy_ddio_dqoe_5,phy_ddio_dqoe_4,phy_ddio_dqoe_3,phy_ddio_dqoe_2,phy_ddio_dqoe_1,phy_ddio_dqoe_0}),
	.write_strobe({phy_ddio_dqs_dout_3,phy_ddio_dqs_dout_2,phy_ddio_dqs_dout_1,phy_ddio_dqs_dout_0}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_0),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_0),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_1,phy_ddio_dqslogic_dqsena_0}),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_1,phy_ddio_dqslogic_dqsena_0}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_0),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_1,phy_ddio_dqslogic_incrdataen_0}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_1,phy_ddio_dqslogic_incwrptr_0}),
	.oct_ena_in({phy_ddio_dqslogic_oct_1,phy_ddio_dqslogic_oct_0}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_4,phy_ddio_dqslogic_readlatency_3,phy_ddio_dqslogic_readlatency_2,phy_ddio_dqslogic_readlatency_1,phy_ddio_dqslogic_readlatency_0}),
	.output_strobe_ena({phy_ddio_dqs_oe_1,phy_ddio_dqs_oe_0}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	config_clock_in,
	hr_clock_in,
	write_strobe_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	lfifo_rdata_en_full,
	vfifo_qvld,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	config_clock_in;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] lfifo_rdata_en_full;
input 	[1:0] vfifo_qvld;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(config_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(config_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_altdqdqs_1 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_4,
	phy_ddio_dmdout_5,
	phy_ddio_dmdout_6,
	phy_ddio_dmdout_7,
	phy_ddio_dqdout_36,
	phy_ddio_dqdout_37,
	phy_ddio_dqdout_38,
	phy_ddio_dqdout_39,
	phy_ddio_dqdout_40,
	phy_ddio_dqdout_41,
	phy_ddio_dqdout_42,
	phy_ddio_dqdout_43,
	phy_ddio_dqdout_44,
	phy_ddio_dqdout_45,
	phy_ddio_dqdout_46,
	phy_ddio_dqdout_47,
	phy_ddio_dqdout_48,
	phy_ddio_dqdout_49,
	phy_ddio_dqdout_50,
	phy_ddio_dqdout_51,
	phy_ddio_dqdout_52,
	phy_ddio_dqdout_53,
	phy_ddio_dqdout_54,
	phy_ddio_dqdout_55,
	phy_ddio_dqdout_56,
	phy_ddio_dqdout_57,
	phy_ddio_dqdout_58,
	phy_ddio_dqdout_59,
	phy_ddio_dqdout_60,
	phy_ddio_dqdout_61,
	phy_ddio_dqdout_62,
	phy_ddio_dqdout_63,
	phy_ddio_dqdout_64,
	phy_ddio_dqdout_65,
	phy_ddio_dqdout_66,
	phy_ddio_dqdout_67,
	phy_ddio_dqoe_18,
	phy_ddio_dqoe_19,
	phy_ddio_dqoe_20,
	phy_ddio_dqoe_21,
	phy_ddio_dqoe_22,
	phy_ddio_dqoe_23,
	phy_ddio_dqoe_24,
	phy_ddio_dqoe_25,
	phy_ddio_dqoe_26,
	phy_ddio_dqoe_27,
	phy_ddio_dqoe_28,
	phy_ddio_dqoe_29,
	phy_ddio_dqoe_30,
	phy_ddio_dqoe_31,
	phy_ddio_dqoe_32,
	phy_ddio_dqoe_33,
	phy_ddio_dqs_dout_4,
	phy_ddio_dqs_dout_5,
	phy_ddio_dqs_dout_6,
	phy_ddio_dqs_dout_7,
	phy_ddio_dqslogic_aclr_fifoctrl_1,
	phy_ddio_dqslogic_aclr_pstamble_1,
	phy_ddio_dqslogic_dqsena_2,
	phy_ddio_dqslogic_dqsena_3,
	phy_ddio_dqslogic_fiforeset_1,
	phy_ddio_dqslogic_incrdataen_2,
	phy_ddio_dqslogic_incrdataen_3,
	phy_ddio_dqslogic_incwrptr_2,
	phy_ddio_dqslogic_incwrptr_3,
	phy_ddio_dqslogic_oct_2,
	phy_ddio_dqslogic_oct_3,
	phy_ddio_dqslogic_readlatency_5,
	phy_ddio_dqslogic_readlatency_6,
	phy_ddio_dqslogic_readlatency_7,
	phy_ddio_dqslogic_readlatency_8,
	phy_ddio_dqslogic_readlatency_9,
	phy_ddio_dqs_oe_2,
	phy_ddio_dqs_oe_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_4;
input 	phy_ddio_dmdout_5;
input 	phy_ddio_dmdout_6;
input 	phy_ddio_dmdout_7;
input 	phy_ddio_dqdout_36;
input 	phy_ddio_dqdout_37;
input 	phy_ddio_dqdout_38;
input 	phy_ddio_dqdout_39;
input 	phy_ddio_dqdout_40;
input 	phy_ddio_dqdout_41;
input 	phy_ddio_dqdout_42;
input 	phy_ddio_dqdout_43;
input 	phy_ddio_dqdout_44;
input 	phy_ddio_dqdout_45;
input 	phy_ddio_dqdout_46;
input 	phy_ddio_dqdout_47;
input 	phy_ddio_dqdout_48;
input 	phy_ddio_dqdout_49;
input 	phy_ddio_dqdout_50;
input 	phy_ddio_dqdout_51;
input 	phy_ddio_dqdout_52;
input 	phy_ddio_dqdout_53;
input 	phy_ddio_dqdout_54;
input 	phy_ddio_dqdout_55;
input 	phy_ddio_dqdout_56;
input 	phy_ddio_dqdout_57;
input 	phy_ddio_dqdout_58;
input 	phy_ddio_dqdout_59;
input 	phy_ddio_dqdout_60;
input 	phy_ddio_dqdout_61;
input 	phy_ddio_dqdout_62;
input 	phy_ddio_dqdout_63;
input 	phy_ddio_dqdout_64;
input 	phy_ddio_dqdout_65;
input 	phy_ddio_dqdout_66;
input 	phy_ddio_dqdout_67;
input 	phy_ddio_dqoe_18;
input 	phy_ddio_dqoe_19;
input 	phy_ddio_dqoe_20;
input 	phy_ddio_dqoe_21;
input 	phy_ddio_dqoe_22;
input 	phy_ddio_dqoe_23;
input 	phy_ddio_dqoe_24;
input 	phy_ddio_dqoe_25;
input 	phy_ddio_dqoe_26;
input 	phy_ddio_dqoe_27;
input 	phy_ddio_dqoe_28;
input 	phy_ddio_dqoe_29;
input 	phy_ddio_dqoe_30;
input 	phy_ddio_dqoe_31;
input 	phy_ddio_dqoe_32;
input 	phy_ddio_dqoe_33;
input 	phy_ddio_dqs_dout_4;
input 	phy_ddio_dqs_dout_5;
input 	phy_ddio_dqs_dout_6;
input 	phy_ddio_dqs_dout_7;
input 	phy_ddio_dqslogic_aclr_fifoctrl_1;
input 	phy_ddio_dqslogic_aclr_pstamble_1;
input 	phy_ddio_dqslogic_dqsena_2;
input 	phy_ddio_dqslogic_dqsena_3;
input 	phy_ddio_dqslogic_fiforeset_1;
input 	phy_ddio_dqslogic_incrdataen_2;
input 	phy_ddio_dqslogic_incrdataen_3;
input 	phy_ddio_dqslogic_incwrptr_2;
input 	phy_ddio_dqslogic_incwrptr_3;
input 	phy_ddio_dqslogic_oct_2;
input 	phy_ddio_dqslogic_oct_3;
input 	phy_ddio_dqslogic_readlatency_5;
input 	phy_ddio_dqslogic_readlatency_6;
input 	phy_ddio_dqslogic_readlatency_7;
input 	phy_ddio_dqslogic_readlatency_8;
input 	phy_ddio_dqslogic_readlatency_9;
input 	phy_ddio_dqs_oe_2;
input 	phy_ddio_dqs_oe_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_1 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.config_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_7,phy_ddio_dmdout_6,phy_ddio_dmdout_5,phy_ddio_dmdout_4}),
	.write_data_in({phy_ddio_dqdout_67,phy_ddio_dqdout_66,phy_ddio_dqdout_65,phy_ddio_dqdout_64,phy_ddio_dqdout_63,phy_ddio_dqdout_62,phy_ddio_dqdout_61,phy_ddio_dqdout_60,phy_ddio_dqdout_59,phy_ddio_dqdout_58,phy_ddio_dqdout_57,phy_ddio_dqdout_56,phy_ddio_dqdout_55,phy_ddio_dqdout_54,
phy_ddio_dqdout_53,phy_ddio_dqdout_52,phy_ddio_dqdout_51,phy_ddio_dqdout_50,phy_ddio_dqdout_49,phy_ddio_dqdout_48,phy_ddio_dqdout_47,phy_ddio_dqdout_46,phy_ddio_dqdout_45,phy_ddio_dqdout_44,phy_ddio_dqdout_43,phy_ddio_dqdout_42,phy_ddio_dqdout_41,phy_ddio_dqdout_40,
phy_ddio_dqdout_39,phy_ddio_dqdout_38,phy_ddio_dqdout_37,phy_ddio_dqdout_36}),
	.write_oe_in({phy_ddio_dqoe_33,phy_ddio_dqoe_32,phy_ddio_dqoe_31,phy_ddio_dqoe_30,phy_ddio_dqoe_29,phy_ddio_dqoe_28,phy_ddio_dqoe_27,phy_ddio_dqoe_26,phy_ddio_dqoe_25,phy_ddio_dqoe_24,phy_ddio_dqoe_23,phy_ddio_dqoe_22,phy_ddio_dqoe_21,phy_ddio_dqoe_20,phy_ddio_dqoe_19,phy_ddio_dqoe_18}),
	.write_strobe({phy_ddio_dqs_dout_7,phy_ddio_dqs_dout_6,phy_ddio_dqs_dout_5,phy_ddio_dqs_dout_4}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_1),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_1),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_3,phy_ddio_dqslogic_dqsena_2}),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_3,phy_ddio_dqslogic_dqsena_2}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_1),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_3,phy_ddio_dqslogic_incrdataen_2}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_3,phy_ddio_dqslogic_incwrptr_2}),
	.oct_ena_in({phy_ddio_dqslogic_oct_3,phy_ddio_dqslogic_oct_2}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_9,phy_ddio_dqslogic_readlatency_8,phy_ddio_dqslogic_readlatency_7,phy_ddio_dqslogic_readlatency_6,phy_ddio_dqslogic_readlatency_5}),
	.output_strobe_ena({phy_ddio_dqs_oe_3,phy_ddio_dqs_oe_2}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_1 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	config_clock_in,
	hr_clock_in,
	write_strobe_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	lfifo_rdata_en_full,
	vfifo_qvld,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	config_clock_in;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] lfifo_rdata_en_full;
input 	[1:0] vfifo_qvld;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(config_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(config_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_altdqdqs_2 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_8,
	phy_ddio_dmdout_9,
	phy_ddio_dmdout_10,
	phy_ddio_dmdout_11,
	phy_ddio_dqdout_72,
	phy_ddio_dqdout_73,
	phy_ddio_dqdout_74,
	phy_ddio_dqdout_75,
	phy_ddio_dqdout_76,
	phy_ddio_dqdout_77,
	phy_ddio_dqdout_78,
	phy_ddio_dqdout_79,
	phy_ddio_dqdout_80,
	phy_ddio_dqdout_81,
	phy_ddio_dqdout_82,
	phy_ddio_dqdout_83,
	phy_ddio_dqdout_84,
	phy_ddio_dqdout_85,
	phy_ddio_dqdout_86,
	phy_ddio_dqdout_87,
	phy_ddio_dqdout_88,
	phy_ddio_dqdout_89,
	phy_ddio_dqdout_90,
	phy_ddio_dqdout_91,
	phy_ddio_dqdout_92,
	phy_ddio_dqdout_93,
	phy_ddio_dqdout_94,
	phy_ddio_dqdout_95,
	phy_ddio_dqdout_96,
	phy_ddio_dqdout_97,
	phy_ddio_dqdout_98,
	phy_ddio_dqdout_99,
	phy_ddio_dqdout_100,
	phy_ddio_dqdout_101,
	phy_ddio_dqdout_102,
	phy_ddio_dqdout_103,
	phy_ddio_dqoe_36,
	phy_ddio_dqoe_37,
	phy_ddio_dqoe_38,
	phy_ddio_dqoe_39,
	phy_ddio_dqoe_40,
	phy_ddio_dqoe_41,
	phy_ddio_dqoe_42,
	phy_ddio_dqoe_43,
	phy_ddio_dqoe_44,
	phy_ddio_dqoe_45,
	phy_ddio_dqoe_46,
	phy_ddio_dqoe_47,
	phy_ddio_dqoe_48,
	phy_ddio_dqoe_49,
	phy_ddio_dqoe_50,
	phy_ddio_dqoe_51,
	phy_ddio_dqs_dout_8,
	phy_ddio_dqs_dout_9,
	phy_ddio_dqs_dout_10,
	phy_ddio_dqs_dout_11,
	phy_ddio_dqslogic_aclr_fifoctrl_2,
	phy_ddio_dqslogic_aclr_pstamble_2,
	phy_ddio_dqslogic_dqsena_4,
	phy_ddio_dqslogic_dqsena_5,
	phy_ddio_dqslogic_fiforeset_2,
	phy_ddio_dqslogic_incrdataen_4,
	phy_ddio_dqslogic_incrdataen_5,
	phy_ddio_dqslogic_incwrptr_4,
	phy_ddio_dqslogic_incwrptr_5,
	phy_ddio_dqslogic_oct_4,
	phy_ddio_dqslogic_oct_5,
	phy_ddio_dqslogic_readlatency_10,
	phy_ddio_dqslogic_readlatency_11,
	phy_ddio_dqslogic_readlatency_12,
	phy_ddio_dqslogic_readlatency_13,
	phy_ddio_dqslogic_readlatency_14,
	phy_ddio_dqs_oe_4,
	phy_ddio_dqs_oe_5,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_8;
input 	phy_ddio_dmdout_9;
input 	phy_ddio_dmdout_10;
input 	phy_ddio_dmdout_11;
input 	phy_ddio_dqdout_72;
input 	phy_ddio_dqdout_73;
input 	phy_ddio_dqdout_74;
input 	phy_ddio_dqdout_75;
input 	phy_ddio_dqdout_76;
input 	phy_ddio_dqdout_77;
input 	phy_ddio_dqdout_78;
input 	phy_ddio_dqdout_79;
input 	phy_ddio_dqdout_80;
input 	phy_ddio_dqdout_81;
input 	phy_ddio_dqdout_82;
input 	phy_ddio_dqdout_83;
input 	phy_ddio_dqdout_84;
input 	phy_ddio_dqdout_85;
input 	phy_ddio_dqdout_86;
input 	phy_ddio_dqdout_87;
input 	phy_ddio_dqdout_88;
input 	phy_ddio_dqdout_89;
input 	phy_ddio_dqdout_90;
input 	phy_ddio_dqdout_91;
input 	phy_ddio_dqdout_92;
input 	phy_ddio_dqdout_93;
input 	phy_ddio_dqdout_94;
input 	phy_ddio_dqdout_95;
input 	phy_ddio_dqdout_96;
input 	phy_ddio_dqdout_97;
input 	phy_ddio_dqdout_98;
input 	phy_ddio_dqdout_99;
input 	phy_ddio_dqdout_100;
input 	phy_ddio_dqdout_101;
input 	phy_ddio_dqdout_102;
input 	phy_ddio_dqdout_103;
input 	phy_ddio_dqoe_36;
input 	phy_ddio_dqoe_37;
input 	phy_ddio_dqoe_38;
input 	phy_ddio_dqoe_39;
input 	phy_ddio_dqoe_40;
input 	phy_ddio_dqoe_41;
input 	phy_ddio_dqoe_42;
input 	phy_ddio_dqoe_43;
input 	phy_ddio_dqoe_44;
input 	phy_ddio_dqoe_45;
input 	phy_ddio_dqoe_46;
input 	phy_ddio_dqoe_47;
input 	phy_ddio_dqoe_48;
input 	phy_ddio_dqoe_49;
input 	phy_ddio_dqoe_50;
input 	phy_ddio_dqoe_51;
input 	phy_ddio_dqs_dout_8;
input 	phy_ddio_dqs_dout_9;
input 	phy_ddio_dqs_dout_10;
input 	phy_ddio_dqs_dout_11;
input 	phy_ddio_dqslogic_aclr_fifoctrl_2;
input 	phy_ddio_dqslogic_aclr_pstamble_2;
input 	phy_ddio_dqslogic_dqsena_4;
input 	phy_ddio_dqslogic_dqsena_5;
input 	phy_ddio_dqslogic_fiforeset_2;
input 	phy_ddio_dqslogic_incrdataen_4;
input 	phy_ddio_dqslogic_incrdataen_5;
input 	phy_ddio_dqslogic_incwrptr_4;
input 	phy_ddio_dqslogic_incwrptr_5;
input 	phy_ddio_dqslogic_oct_4;
input 	phy_ddio_dqslogic_oct_5;
input 	phy_ddio_dqslogic_readlatency_10;
input 	phy_ddio_dqslogic_readlatency_11;
input 	phy_ddio_dqslogic_readlatency_12;
input 	phy_ddio_dqslogic_readlatency_13;
input 	phy_ddio_dqslogic_readlatency_14;
input 	phy_ddio_dqs_oe_4;
input 	phy_ddio_dqs_oe_5;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_2 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.config_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_11,phy_ddio_dmdout_10,phy_ddio_dmdout_9,phy_ddio_dmdout_8}),
	.write_data_in({phy_ddio_dqdout_103,phy_ddio_dqdout_102,phy_ddio_dqdout_101,phy_ddio_dqdout_100,phy_ddio_dqdout_99,phy_ddio_dqdout_98,phy_ddio_dqdout_97,phy_ddio_dqdout_96,phy_ddio_dqdout_95,phy_ddio_dqdout_94,phy_ddio_dqdout_93,phy_ddio_dqdout_92,phy_ddio_dqdout_91,phy_ddio_dqdout_90,
phy_ddio_dqdout_89,phy_ddio_dqdout_88,phy_ddio_dqdout_87,phy_ddio_dqdout_86,phy_ddio_dqdout_85,phy_ddio_dqdout_84,phy_ddio_dqdout_83,phy_ddio_dqdout_82,phy_ddio_dqdout_81,phy_ddio_dqdout_80,phy_ddio_dqdout_79,phy_ddio_dqdout_78,phy_ddio_dqdout_77,phy_ddio_dqdout_76,
phy_ddio_dqdout_75,phy_ddio_dqdout_74,phy_ddio_dqdout_73,phy_ddio_dqdout_72}),
	.write_oe_in({phy_ddio_dqoe_51,phy_ddio_dqoe_50,phy_ddio_dqoe_49,phy_ddio_dqoe_48,phy_ddio_dqoe_47,phy_ddio_dqoe_46,phy_ddio_dqoe_45,phy_ddio_dqoe_44,phy_ddio_dqoe_43,phy_ddio_dqoe_42,phy_ddio_dqoe_41,phy_ddio_dqoe_40,phy_ddio_dqoe_39,phy_ddio_dqoe_38,phy_ddio_dqoe_37,phy_ddio_dqoe_36}),
	.write_strobe({phy_ddio_dqs_dout_11,phy_ddio_dqs_dout_10,phy_ddio_dqs_dout_9,phy_ddio_dqs_dout_8}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_2),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_2),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_5,phy_ddio_dqslogic_dqsena_4}),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_5,phy_ddio_dqslogic_dqsena_4}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_2),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_5,phy_ddio_dqslogic_incrdataen_4}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_5,phy_ddio_dqslogic_incwrptr_4}),
	.oct_ena_in({phy_ddio_dqslogic_oct_5,phy_ddio_dqslogic_oct_4}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_14,phy_ddio_dqslogic_readlatency_13,phy_ddio_dqslogic_readlatency_12,phy_ddio_dqslogic_readlatency_11,phy_ddio_dqslogic_readlatency_10}),
	.output_strobe_ena({phy_ddio_dqs_oe_5,phy_ddio_dqs_oe_4}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_2 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	config_clock_in,
	hr_clock_in,
	write_strobe_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	lfifo_rdata_en_full,
	vfifo_qvld,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	config_clock_in;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] lfifo_rdata_en_full;
input 	[1:0] vfifo_qvld;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(config_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(config_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_altdqdqs_3 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_12,
	phy_ddio_dmdout_13,
	phy_ddio_dmdout_14,
	phy_ddio_dmdout_15,
	phy_ddio_dqdout_108,
	phy_ddio_dqdout_109,
	phy_ddio_dqdout_110,
	phy_ddio_dqdout_111,
	phy_ddio_dqdout_112,
	phy_ddio_dqdout_113,
	phy_ddio_dqdout_114,
	phy_ddio_dqdout_115,
	phy_ddio_dqdout_116,
	phy_ddio_dqdout_117,
	phy_ddio_dqdout_118,
	phy_ddio_dqdout_119,
	phy_ddio_dqdout_120,
	phy_ddio_dqdout_121,
	phy_ddio_dqdout_122,
	phy_ddio_dqdout_123,
	phy_ddio_dqdout_124,
	phy_ddio_dqdout_125,
	phy_ddio_dqdout_126,
	phy_ddio_dqdout_127,
	phy_ddio_dqdout_128,
	phy_ddio_dqdout_129,
	phy_ddio_dqdout_130,
	phy_ddio_dqdout_131,
	phy_ddio_dqdout_132,
	phy_ddio_dqdout_133,
	phy_ddio_dqdout_134,
	phy_ddio_dqdout_135,
	phy_ddio_dqdout_136,
	phy_ddio_dqdout_137,
	phy_ddio_dqdout_138,
	phy_ddio_dqdout_139,
	phy_ddio_dqoe_54,
	phy_ddio_dqoe_55,
	phy_ddio_dqoe_56,
	phy_ddio_dqoe_57,
	phy_ddio_dqoe_58,
	phy_ddio_dqoe_59,
	phy_ddio_dqoe_60,
	phy_ddio_dqoe_61,
	phy_ddio_dqoe_62,
	phy_ddio_dqoe_63,
	phy_ddio_dqoe_64,
	phy_ddio_dqoe_65,
	phy_ddio_dqoe_66,
	phy_ddio_dqoe_67,
	phy_ddio_dqoe_68,
	phy_ddio_dqoe_69,
	phy_ddio_dqs_dout_12,
	phy_ddio_dqs_dout_13,
	phy_ddio_dqs_dout_14,
	phy_ddio_dqs_dout_15,
	phy_ddio_dqslogic_aclr_fifoctrl_3,
	phy_ddio_dqslogic_aclr_pstamble_3,
	phy_ddio_dqslogic_dqsena_6,
	phy_ddio_dqslogic_dqsena_7,
	phy_ddio_dqslogic_fiforeset_3,
	phy_ddio_dqslogic_incrdataen_6,
	phy_ddio_dqslogic_incrdataen_7,
	phy_ddio_dqslogic_incwrptr_6,
	phy_ddio_dqslogic_incwrptr_7,
	phy_ddio_dqslogic_oct_6,
	phy_ddio_dqslogic_oct_7,
	phy_ddio_dqslogic_readlatency_15,
	phy_ddio_dqslogic_readlatency_16,
	phy_ddio_dqslogic_readlatency_17,
	phy_ddio_dqslogic_readlatency_18,
	phy_ddio_dqslogic_readlatency_19,
	phy_ddio_dqs_oe_6,
	phy_ddio_dqs_oe_7,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_12;
input 	phy_ddio_dmdout_13;
input 	phy_ddio_dmdout_14;
input 	phy_ddio_dmdout_15;
input 	phy_ddio_dqdout_108;
input 	phy_ddio_dqdout_109;
input 	phy_ddio_dqdout_110;
input 	phy_ddio_dqdout_111;
input 	phy_ddio_dqdout_112;
input 	phy_ddio_dqdout_113;
input 	phy_ddio_dqdout_114;
input 	phy_ddio_dqdout_115;
input 	phy_ddio_dqdout_116;
input 	phy_ddio_dqdout_117;
input 	phy_ddio_dqdout_118;
input 	phy_ddio_dqdout_119;
input 	phy_ddio_dqdout_120;
input 	phy_ddio_dqdout_121;
input 	phy_ddio_dqdout_122;
input 	phy_ddio_dqdout_123;
input 	phy_ddio_dqdout_124;
input 	phy_ddio_dqdout_125;
input 	phy_ddio_dqdout_126;
input 	phy_ddio_dqdout_127;
input 	phy_ddio_dqdout_128;
input 	phy_ddio_dqdout_129;
input 	phy_ddio_dqdout_130;
input 	phy_ddio_dqdout_131;
input 	phy_ddio_dqdout_132;
input 	phy_ddio_dqdout_133;
input 	phy_ddio_dqdout_134;
input 	phy_ddio_dqdout_135;
input 	phy_ddio_dqdout_136;
input 	phy_ddio_dqdout_137;
input 	phy_ddio_dqdout_138;
input 	phy_ddio_dqdout_139;
input 	phy_ddio_dqoe_54;
input 	phy_ddio_dqoe_55;
input 	phy_ddio_dqoe_56;
input 	phy_ddio_dqoe_57;
input 	phy_ddio_dqoe_58;
input 	phy_ddio_dqoe_59;
input 	phy_ddio_dqoe_60;
input 	phy_ddio_dqoe_61;
input 	phy_ddio_dqoe_62;
input 	phy_ddio_dqoe_63;
input 	phy_ddio_dqoe_64;
input 	phy_ddio_dqoe_65;
input 	phy_ddio_dqoe_66;
input 	phy_ddio_dqoe_67;
input 	phy_ddio_dqoe_68;
input 	phy_ddio_dqoe_69;
input 	phy_ddio_dqs_dout_12;
input 	phy_ddio_dqs_dout_13;
input 	phy_ddio_dqs_dout_14;
input 	phy_ddio_dqs_dout_15;
input 	phy_ddio_dqslogic_aclr_fifoctrl_3;
input 	phy_ddio_dqslogic_aclr_pstamble_3;
input 	phy_ddio_dqslogic_dqsena_6;
input 	phy_ddio_dqslogic_dqsena_7;
input 	phy_ddio_dqslogic_fiforeset_3;
input 	phy_ddio_dqslogic_incrdataen_6;
input 	phy_ddio_dqslogic_incrdataen_7;
input 	phy_ddio_dqslogic_incwrptr_6;
input 	phy_ddio_dqslogic_incwrptr_7;
input 	phy_ddio_dqslogic_oct_6;
input 	phy_ddio_dqslogic_oct_7;
input 	phy_ddio_dqslogic_readlatency_15;
input 	phy_ddio_dqslogic_readlatency_16;
input 	phy_ddio_dqslogic_readlatency_17;
input 	phy_ddio_dqslogic_readlatency_18;
input 	phy_ddio_dqslogic_readlatency_19;
input 	phy_ddio_dqs_oe_6;
input 	phy_ddio_dqs_oe_7;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_3 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.config_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_15,phy_ddio_dmdout_14,phy_ddio_dmdout_13,phy_ddio_dmdout_12}),
	.write_data_in({phy_ddio_dqdout_139,phy_ddio_dqdout_138,phy_ddio_dqdout_137,phy_ddio_dqdout_136,phy_ddio_dqdout_135,phy_ddio_dqdout_134,phy_ddio_dqdout_133,phy_ddio_dqdout_132,phy_ddio_dqdout_131,phy_ddio_dqdout_130,phy_ddio_dqdout_129,phy_ddio_dqdout_128,phy_ddio_dqdout_127,
phy_ddio_dqdout_126,phy_ddio_dqdout_125,phy_ddio_dqdout_124,phy_ddio_dqdout_123,phy_ddio_dqdout_122,phy_ddio_dqdout_121,phy_ddio_dqdout_120,phy_ddio_dqdout_119,phy_ddio_dqdout_118,phy_ddio_dqdout_117,phy_ddio_dqdout_116,phy_ddio_dqdout_115,phy_ddio_dqdout_114,
phy_ddio_dqdout_113,phy_ddio_dqdout_112,phy_ddio_dqdout_111,phy_ddio_dqdout_110,phy_ddio_dqdout_109,phy_ddio_dqdout_108}),
	.write_oe_in({phy_ddio_dqoe_69,phy_ddio_dqoe_68,phy_ddio_dqoe_67,phy_ddio_dqoe_66,phy_ddio_dqoe_65,phy_ddio_dqoe_64,phy_ddio_dqoe_63,phy_ddio_dqoe_62,phy_ddio_dqoe_61,phy_ddio_dqoe_60,phy_ddio_dqoe_59,phy_ddio_dqoe_58,phy_ddio_dqoe_57,phy_ddio_dqoe_56,phy_ddio_dqoe_55,phy_ddio_dqoe_54}),
	.write_strobe({phy_ddio_dqs_dout_15,phy_ddio_dqs_dout_14,phy_ddio_dqs_dout_13,phy_ddio_dqs_dout_12}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_3),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_3),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_7,phy_ddio_dqslogic_dqsena_6}),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_7,phy_ddio_dqslogic_dqsena_6}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_3),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_7,phy_ddio_dqslogic_incrdataen_6}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_7,phy_ddio_dqslogic_incwrptr_6}),
	.oct_ena_in({phy_ddio_dqslogic_oct_7,phy_ddio_dqslogic_oct_6}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_19,phy_ddio_dqslogic_readlatency_18,phy_ddio_dqslogic_readlatency_17,phy_ddio_dqslogic_readlatency_16,phy_ddio_dqslogic_readlatency_15}),
	.output_strobe_ena({phy_ddio_dqs_oe_7,phy_ddio_dqs_oe_6}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module Computer_System_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_3 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	config_clock_in,
	hr_clock_in,
	write_strobe_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	lfifo_rdata_en_full,
	vfifo_qvld,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	config_clock_in;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] lfifo_rdata_en_full;
input 	[1:0] vfifo_qvld;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(config_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(config_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module Computer_System_hps_sdram_p0_acv_ldc_25 (
	pll_dqs_clk,
	pll_hr_clk,
	afi_clk,
	avl_clk,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
input 	pll_hr_clk;
output 	afi_clk;
output 	avl_clk;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;

assign afi_clk = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

assign avl_clk = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(pll_dqs_clk),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

endmodule

module Computer_System_hps_sdram_pll (
	pll_mem_clk,
	pll_write_clk)/* synthesis synthesis_greybox=0 */;
output 	pll_mem_clk;
output 	pll_write_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \clk_out[2] ;
wire \clk_out[3] ;

wire [3:0] pll_CLK_OUT_bus;

assign pll_mem_clk = pll_CLK_OUT_bus[0];
assign pll_write_clk = pll_CLK_OUT_bus[1];
assign \clk_out[2]  = pll_CLK_OUT_bus[2];
assign \clk_out[3]  = pll_CLK_OUT_bus[3];

cyclonev_hps_sdram_pll pll(
	.ref_clk(gnd),
	.clk_out(pll_CLK_OUT_bus));

endmodule

module Computer_System_Computer_System_fifo_HPS_to_FPGA (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	outclk_wire_0,
	op_2,
	op_21,
	op_22,
	aneb_result_wire_0,
	rdclk_control_slave_readdata_0,
	rdclk_control_slave_readdata_1,
	rdclk_control_slave_readdata_2,
	rdclk_control_slave_readdata_3,
	rdclk_control_slave_readdata_4,
	rdclk_control_slave_readdata_5,
	rdclk_control_slave_readdata_6,
	rdclk_control_slave_readdata_7,
	wait_latency_counter_0,
	wait_latency_counter_1,
	avalonmm_write_slave_waitrequest,
	wrfull,
	wrfull1,
	m0_write,
	in_data_reg_0,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	r_sync_rst,
	r_sync_rst1,
	m0_write1,
	m0_read,
	wrclk_control_slave_readdata_0,
	wrclk_control_slave_readdata_1,
	wrclk_control_slave_readdata_2,
	wrclk_control_slave_readdata_3,
	wrclk_control_slave_readdata_4,
	wrclk_control_slave_readdata_5,
	wrclk_control_slave_readdata_6,
	wrclk_control_slave_readdata_7,
	wrfull2,
	wrfull3,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_3,
	in_data_reg_01,
	in_data_reg_210,
	in_data_reg_110,
	in_data_reg_141,
	in_data_reg_81,
	in_data_reg_131,
	in_data_reg_121,
	in_data_reg_111,
	in_data_reg_101,
	in_data_reg_91,
	in_data_reg_191,
	in_data_reg_181,
	in_data_reg_171,
	in_data_reg_161,
	in_data_reg_151,
	in_data_reg_261,
	in_data_reg_211,
	in_data_reg_201,
	in_data_reg_311,
	in_data_reg_301,
	in_data_reg_291,
	in_data_reg_281,
	in_data_reg_271,
	in_data_reg_251,
	in_data_reg_241,
	in_data_reg_231,
	in_data_reg_221,
	in_data_reg_71,
	in_data_reg_61,
	in_data_reg_51,
	in_data_reg_41,
	in_data_reg_32,
	fifo_hps_to_fpga_out_read,
	clock_bridge_0_in_clk_clk,
	fifo_hps_to_fpga_out_csr_address_2,
	fifo_hps_to_fpga_out_csr_address_0,
	fifo_hps_to_fpga_out_csr_address_1,
	fifo_hps_to_fpga_out_csr_read,
	fifo_hps_to_fpga_out_csr_writedata_0,
	fifo_hps_to_fpga_out_csr_write,
	fifo_hps_to_fpga_out_csr_writedata_7,
	fifo_hps_to_fpga_out_csr_writedata_1,
	fifo_hps_to_fpga_out_csr_writedata_13,
	fifo_hps_to_fpga_out_csr_writedata_19,
	fifo_hps_to_fpga_out_csr_writedata_26,
	fifo_hps_to_fpga_out_csr_writedata_27,
	fifo_hps_to_fpga_out_csr_writedata_28,
	fifo_hps_to_fpga_out_csr_writedata_29,
	fifo_hps_to_fpga_out_csr_writedata_30,
	fifo_hps_to_fpga_out_csr_writedata_31,
	fifo_hps_to_fpga_out_csr_writedata_20,
	fifo_hps_to_fpga_out_csr_writedata_21,
	fifo_hps_to_fpga_out_csr_writedata_22,
	fifo_hps_to_fpga_out_csr_writedata_23,
	fifo_hps_to_fpga_out_csr_writedata_24,
	fifo_hps_to_fpga_out_csr_writedata_25,
	fifo_hps_to_fpga_out_csr_writedata_8,
	fifo_hps_to_fpga_out_csr_writedata_9,
	fifo_hps_to_fpga_out_csr_writedata_10,
	fifo_hps_to_fpga_out_csr_writedata_11,
	fifo_hps_to_fpga_out_csr_writedata_12,
	fifo_hps_to_fpga_out_csr_writedata_14,
	fifo_hps_to_fpga_out_csr_writedata_15,
	fifo_hps_to_fpga_out_csr_writedata_16,
	fifo_hps_to_fpga_out_csr_writedata_17,
	fifo_hps_to_fpga_out_csr_writedata_18,
	fifo_hps_to_fpga_out_csr_writedata_2,
	fifo_hps_to_fpga_out_csr_writedata_3,
	fifo_hps_to_fpga_out_csr_writedata_4,
	fifo_hps_to_fpga_out_csr_writedata_5,
	fifo_hps_to_fpga_out_csr_writedata_6)/* synthesis synthesis_greybox=0 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
input 	outclk_wire_0;
output 	op_2;
output 	op_21;
output 	op_22;
output 	aneb_result_wire_0;
output 	rdclk_control_slave_readdata_0;
output 	rdclk_control_slave_readdata_1;
output 	rdclk_control_slave_readdata_2;
output 	rdclk_control_slave_readdata_3;
output 	rdclk_control_slave_readdata_4;
output 	rdclk_control_slave_readdata_5;
output 	rdclk_control_slave_readdata_6;
output 	rdclk_control_slave_readdata_7;
input 	wait_latency_counter_0;
input 	wait_latency_counter_1;
output 	avalonmm_write_slave_waitrequest;
output 	wrfull;
output 	wrfull1;
input 	m0_write;
input 	in_data_reg_0;
input 	in_data_reg_1;
input 	in_data_reg_2;
input 	in_data_reg_3;
input 	in_data_reg_4;
input 	in_data_reg_5;
input 	in_data_reg_6;
input 	in_data_reg_7;
input 	in_data_reg_8;
input 	in_data_reg_9;
input 	in_data_reg_10;
input 	in_data_reg_11;
input 	in_data_reg_12;
input 	in_data_reg_13;
input 	in_data_reg_14;
input 	in_data_reg_15;
input 	in_data_reg_16;
input 	in_data_reg_17;
input 	in_data_reg_18;
input 	in_data_reg_19;
input 	in_data_reg_20;
input 	in_data_reg_21;
input 	in_data_reg_22;
input 	in_data_reg_23;
input 	in_data_reg_24;
input 	in_data_reg_25;
input 	in_data_reg_26;
input 	in_data_reg_27;
input 	in_data_reg_28;
input 	in_data_reg_29;
input 	in_data_reg_30;
input 	in_data_reg_31;
input 	r_sync_rst;
input 	r_sync_rst1;
input 	m0_write1;
input 	m0_read;
output 	wrclk_control_slave_readdata_0;
output 	wrclk_control_slave_readdata_1;
output 	wrclk_control_slave_readdata_2;
output 	wrclk_control_slave_readdata_3;
output 	wrclk_control_slave_readdata_4;
output 	wrclk_control_slave_readdata_5;
output 	wrclk_control_slave_readdata_6;
output 	wrclk_control_slave_readdata_7;
output 	wrfull2;
output 	wrfull3;
input 	int_nxt_addr_reg_dly_2;
input 	int_nxt_addr_reg_dly_4;
input 	int_nxt_addr_reg_dly_3;
input 	in_data_reg_01;
input 	in_data_reg_210;
input 	in_data_reg_110;
input 	in_data_reg_141;
input 	in_data_reg_81;
input 	in_data_reg_131;
input 	in_data_reg_121;
input 	in_data_reg_111;
input 	in_data_reg_101;
input 	in_data_reg_91;
input 	in_data_reg_191;
input 	in_data_reg_181;
input 	in_data_reg_171;
input 	in_data_reg_161;
input 	in_data_reg_151;
input 	in_data_reg_261;
input 	in_data_reg_211;
input 	in_data_reg_201;
input 	in_data_reg_311;
input 	in_data_reg_301;
input 	in_data_reg_291;
input 	in_data_reg_281;
input 	in_data_reg_271;
input 	in_data_reg_251;
input 	in_data_reg_241;
input 	in_data_reg_231;
input 	in_data_reg_221;
input 	in_data_reg_71;
input 	in_data_reg_61;
input 	in_data_reg_51;
input 	in_data_reg_41;
input 	in_data_reg_32;
input 	fifo_hps_to_fpga_out_read;
input 	clock_bridge_0_in_clk_clk;
input 	fifo_hps_to_fpga_out_csr_address_2;
input 	fifo_hps_to_fpga_out_csr_address_0;
input 	fifo_hps_to_fpga_out_csr_address_1;
input 	fifo_hps_to_fpga_out_csr_read;
input 	fifo_hps_to_fpga_out_csr_writedata_0;
input 	fifo_hps_to_fpga_out_csr_write;
input 	fifo_hps_to_fpga_out_csr_writedata_7;
input 	fifo_hps_to_fpga_out_csr_writedata_1;
input 	fifo_hps_to_fpga_out_csr_writedata_13;
input 	fifo_hps_to_fpga_out_csr_writedata_19;
input 	fifo_hps_to_fpga_out_csr_writedata_26;
input 	fifo_hps_to_fpga_out_csr_writedata_27;
input 	fifo_hps_to_fpga_out_csr_writedata_28;
input 	fifo_hps_to_fpga_out_csr_writedata_29;
input 	fifo_hps_to_fpga_out_csr_writedata_30;
input 	fifo_hps_to_fpga_out_csr_writedata_31;
input 	fifo_hps_to_fpga_out_csr_writedata_20;
input 	fifo_hps_to_fpga_out_csr_writedata_21;
input 	fifo_hps_to_fpga_out_csr_writedata_22;
input 	fifo_hps_to_fpga_out_csr_writedata_23;
input 	fifo_hps_to_fpga_out_csr_writedata_24;
input 	fifo_hps_to_fpga_out_csr_writedata_25;
input 	fifo_hps_to_fpga_out_csr_writedata_8;
input 	fifo_hps_to_fpga_out_csr_writedata_9;
input 	fifo_hps_to_fpga_out_csr_writedata_10;
input 	fifo_hps_to_fpga_out_csr_writedata_11;
input 	fifo_hps_to_fpga_out_csr_writedata_12;
input 	fifo_hps_to_fpga_out_csr_writedata_14;
input 	fifo_hps_to_fpga_out_csr_writedata_15;
input 	fifo_hps_to_fpga_out_csr_writedata_16;
input 	fifo_hps_to_fpga_out_csr_writedata_17;
input 	fifo_hps_to_fpga_out_csr_writedata_18;
input 	fifo_hps_to_fpga_out_csr_writedata_2;
input 	fifo_hps_to_fpga_out_csr_writedata_3;
input 	fifo_hps_to_fpga_out_csr_writedata_4;
input 	fifo_hps_to_fpga_out_csr_writedata_5;
input 	fifo_hps_to_fpga_out_csr_writedata_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls the_dcfifo_with_controls(
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.outclk_wire_0(outclk_wire_0),
	.op_2(op_2),
	.op_21(op_21),
	.op_22(op_22),
	.aneb_result_wire_0(aneb_result_wire_0),
	.rdclk_control_slave_readdata_0(rdclk_control_slave_readdata_0),
	.rdclk_control_slave_readdata_1(rdclk_control_slave_readdata_1),
	.rdclk_control_slave_readdata_2(rdclk_control_slave_readdata_2),
	.rdclk_control_slave_readdata_3(rdclk_control_slave_readdata_3),
	.rdclk_control_slave_readdata_4(rdclk_control_slave_readdata_4),
	.rdclk_control_slave_readdata_5(rdclk_control_slave_readdata_5),
	.rdclk_control_slave_readdata_6(rdclk_control_slave_readdata_6),
	.rdclk_control_slave_readdata_7(rdclk_control_slave_readdata_7),
	.wait_latency_counter_0(wait_latency_counter_0),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wrfull(avalonmm_write_slave_waitrequest),
	.wrfull1(wrfull),
	.wrfull2(wrfull1),
	.m0_write(m0_write),
	.in_data_reg_0(in_data_reg_0),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_24(in_data_reg_24),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_31(in_data_reg_31),
	.r_sync_rst(r_sync_rst),
	.r_sync_rst1(r_sync_rst1),
	.m0_write1(m0_write1),
	.m0_read(m0_read),
	.wrclk_control_slave_readdata_0(wrclk_control_slave_readdata_0),
	.wrclk_control_slave_readdata_1(wrclk_control_slave_readdata_1),
	.wrclk_control_slave_readdata_2(wrclk_control_slave_readdata_2),
	.wrclk_control_slave_readdata_3(wrclk_control_slave_readdata_3),
	.wrclk_control_slave_readdata_4(wrclk_control_slave_readdata_4),
	.wrclk_control_slave_readdata_5(wrclk_control_slave_readdata_5),
	.wrclk_control_slave_readdata_6(wrclk_control_slave_readdata_6),
	.wrclk_control_slave_readdata_7(wrclk_control_slave_readdata_7),
	.wrfull3(wrfull2),
	.wrfull4(wrfull3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_4(int_nxt_addr_reg_dly_4),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.wrclk_control_slave_writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,in_data_reg_51,in_data_reg_41,in_data_reg_32,in_data_reg_210,in_data_reg_110,in_data_reg_01}),
	.in_data_reg_141(in_data_reg_141),
	.in_data_reg_81(in_data_reg_81),
	.in_data_reg_131(in_data_reg_131),
	.in_data_reg_121(in_data_reg_121),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_101(in_data_reg_101),
	.in_data_reg_91(in_data_reg_91),
	.in_data_reg_191(in_data_reg_191),
	.in_data_reg_181(in_data_reg_181),
	.in_data_reg_171(in_data_reg_171),
	.in_data_reg_161(in_data_reg_161),
	.in_data_reg_151(in_data_reg_151),
	.in_data_reg_261(in_data_reg_261),
	.in_data_reg_211(in_data_reg_211),
	.in_data_reg_201(in_data_reg_201),
	.in_data_reg_311(in_data_reg_311),
	.in_data_reg_301(in_data_reg_301),
	.in_data_reg_291(in_data_reg_291),
	.in_data_reg_281(in_data_reg_281),
	.in_data_reg_271(in_data_reg_271),
	.in_data_reg_251(in_data_reg_251),
	.in_data_reg_241(in_data_reg_241),
	.in_data_reg_231(in_data_reg_231),
	.in_data_reg_221(in_data_reg_221),
	.in_data_reg_71(in_data_reg_71),
	.in_data_reg_61(in_data_reg_61),
	.fifo_hps_to_fpga_out_read(fifo_hps_to_fpga_out_read),
	.clock_bridge_0_in_clk_clk(clock_bridge_0_in_clk_clk),
	.fifo_hps_to_fpga_out_csr_address_2(fifo_hps_to_fpga_out_csr_address_2),
	.fifo_hps_to_fpga_out_csr_address_0(fifo_hps_to_fpga_out_csr_address_0),
	.fifo_hps_to_fpga_out_csr_address_1(fifo_hps_to_fpga_out_csr_address_1),
	.fifo_hps_to_fpga_out_csr_read(fifo_hps_to_fpga_out_csr_read),
	.rdclk_control_slave_writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,fifo_hps_to_fpga_out_csr_writedata_5,fifo_hps_to_fpga_out_csr_writedata_4,fifo_hps_to_fpga_out_csr_writedata_3,fifo_hps_to_fpga_out_csr_writedata_2,
fifo_hps_to_fpga_out_csr_writedata_1,fifo_hps_to_fpga_out_csr_writedata_0}),
	.fifo_hps_to_fpga_out_csr_write(fifo_hps_to_fpga_out_csr_write),
	.fifo_hps_to_fpga_out_csr_writedata_7(fifo_hps_to_fpga_out_csr_writedata_7),
	.fifo_hps_to_fpga_out_csr_writedata_13(fifo_hps_to_fpga_out_csr_writedata_13),
	.fifo_hps_to_fpga_out_csr_writedata_19(fifo_hps_to_fpga_out_csr_writedata_19),
	.fifo_hps_to_fpga_out_csr_writedata_26(fifo_hps_to_fpga_out_csr_writedata_26),
	.fifo_hps_to_fpga_out_csr_writedata_27(fifo_hps_to_fpga_out_csr_writedata_27),
	.fifo_hps_to_fpga_out_csr_writedata_28(fifo_hps_to_fpga_out_csr_writedata_28),
	.fifo_hps_to_fpga_out_csr_writedata_29(fifo_hps_to_fpga_out_csr_writedata_29),
	.fifo_hps_to_fpga_out_csr_writedata_30(fifo_hps_to_fpga_out_csr_writedata_30),
	.fifo_hps_to_fpga_out_csr_writedata_31(fifo_hps_to_fpga_out_csr_writedata_31),
	.fifo_hps_to_fpga_out_csr_writedata_20(fifo_hps_to_fpga_out_csr_writedata_20),
	.fifo_hps_to_fpga_out_csr_writedata_21(fifo_hps_to_fpga_out_csr_writedata_21),
	.fifo_hps_to_fpga_out_csr_writedata_22(fifo_hps_to_fpga_out_csr_writedata_22),
	.fifo_hps_to_fpga_out_csr_writedata_23(fifo_hps_to_fpga_out_csr_writedata_23),
	.fifo_hps_to_fpga_out_csr_writedata_24(fifo_hps_to_fpga_out_csr_writedata_24),
	.fifo_hps_to_fpga_out_csr_writedata_25(fifo_hps_to_fpga_out_csr_writedata_25),
	.fifo_hps_to_fpga_out_csr_writedata_8(fifo_hps_to_fpga_out_csr_writedata_8),
	.fifo_hps_to_fpga_out_csr_writedata_9(fifo_hps_to_fpga_out_csr_writedata_9),
	.fifo_hps_to_fpga_out_csr_writedata_10(fifo_hps_to_fpga_out_csr_writedata_10),
	.fifo_hps_to_fpga_out_csr_writedata_11(fifo_hps_to_fpga_out_csr_writedata_11),
	.fifo_hps_to_fpga_out_csr_writedata_12(fifo_hps_to_fpga_out_csr_writedata_12),
	.fifo_hps_to_fpga_out_csr_writedata_14(fifo_hps_to_fpga_out_csr_writedata_14),
	.fifo_hps_to_fpga_out_csr_writedata_15(fifo_hps_to_fpga_out_csr_writedata_15),
	.fifo_hps_to_fpga_out_csr_writedata_16(fifo_hps_to_fpga_out_csr_writedata_16),
	.fifo_hps_to_fpga_out_csr_writedata_17(fifo_hps_to_fpga_out_csr_writedata_17),
	.fifo_hps_to_fpga_out_csr_writedata_18(fifo_hps_to_fpga_out_csr_writedata_18),
	.fifo_hps_to_fpga_out_csr_writedata_6(fifo_hps_to_fpga_out_csr_writedata_6));

endmodule

module Computer_System_Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	outclk_wire_0,
	op_2,
	op_21,
	op_22,
	aneb_result_wire_0,
	rdclk_control_slave_readdata_0,
	rdclk_control_slave_readdata_1,
	rdclk_control_slave_readdata_2,
	rdclk_control_slave_readdata_3,
	rdclk_control_slave_readdata_4,
	rdclk_control_slave_readdata_5,
	rdclk_control_slave_readdata_6,
	rdclk_control_slave_readdata_7,
	wait_latency_counter_0,
	wait_latency_counter_1,
	wrfull,
	wrfull1,
	wrfull2,
	m0_write,
	in_data_reg_0,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	r_sync_rst,
	r_sync_rst1,
	m0_write1,
	m0_read,
	wrclk_control_slave_readdata_0,
	wrclk_control_slave_readdata_1,
	wrclk_control_slave_readdata_2,
	wrclk_control_slave_readdata_3,
	wrclk_control_slave_readdata_4,
	wrclk_control_slave_readdata_5,
	wrclk_control_slave_readdata_6,
	wrclk_control_slave_readdata_7,
	wrfull3,
	wrfull4,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_3,
	wrclk_control_slave_writedata,
	in_data_reg_141,
	in_data_reg_81,
	in_data_reg_131,
	in_data_reg_121,
	in_data_reg_111,
	in_data_reg_101,
	in_data_reg_91,
	in_data_reg_191,
	in_data_reg_181,
	in_data_reg_171,
	in_data_reg_161,
	in_data_reg_151,
	in_data_reg_261,
	in_data_reg_211,
	in_data_reg_201,
	in_data_reg_311,
	in_data_reg_301,
	in_data_reg_291,
	in_data_reg_281,
	in_data_reg_271,
	in_data_reg_251,
	in_data_reg_241,
	in_data_reg_231,
	in_data_reg_221,
	in_data_reg_71,
	in_data_reg_61,
	fifo_hps_to_fpga_out_read,
	clock_bridge_0_in_clk_clk,
	fifo_hps_to_fpga_out_csr_address_2,
	fifo_hps_to_fpga_out_csr_address_0,
	fifo_hps_to_fpga_out_csr_address_1,
	fifo_hps_to_fpga_out_csr_read,
	rdclk_control_slave_writedata,
	fifo_hps_to_fpga_out_csr_write,
	fifo_hps_to_fpga_out_csr_writedata_7,
	fifo_hps_to_fpga_out_csr_writedata_13,
	fifo_hps_to_fpga_out_csr_writedata_19,
	fifo_hps_to_fpga_out_csr_writedata_26,
	fifo_hps_to_fpga_out_csr_writedata_27,
	fifo_hps_to_fpga_out_csr_writedata_28,
	fifo_hps_to_fpga_out_csr_writedata_29,
	fifo_hps_to_fpga_out_csr_writedata_30,
	fifo_hps_to_fpga_out_csr_writedata_31,
	fifo_hps_to_fpga_out_csr_writedata_20,
	fifo_hps_to_fpga_out_csr_writedata_21,
	fifo_hps_to_fpga_out_csr_writedata_22,
	fifo_hps_to_fpga_out_csr_writedata_23,
	fifo_hps_to_fpga_out_csr_writedata_24,
	fifo_hps_to_fpga_out_csr_writedata_25,
	fifo_hps_to_fpga_out_csr_writedata_8,
	fifo_hps_to_fpga_out_csr_writedata_9,
	fifo_hps_to_fpga_out_csr_writedata_10,
	fifo_hps_to_fpga_out_csr_writedata_11,
	fifo_hps_to_fpga_out_csr_writedata_12,
	fifo_hps_to_fpga_out_csr_writedata_14,
	fifo_hps_to_fpga_out_csr_writedata_15,
	fifo_hps_to_fpga_out_csr_writedata_16,
	fifo_hps_to_fpga_out_csr_writedata_17,
	fifo_hps_to_fpga_out_csr_writedata_18,
	fifo_hps_to_fpga_out_csr_writedata_6)/* synthesis synthesis_greybox=0 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
input 	outclk_wire_0;
output 	op_2;
output 	op_21;
output 	op_22;
output 	aneb_result_wire_0;
output 	rdclk_control_slave_readdata_0;
output 	rdclk_control_slave_readdata_1;
output 	rdclk_control_slave_readdata_2;
output 	rdclk_control_slave_readdata_3;
output 	rdclk_control_slave_readdata_4;
output 	rdclk_control_slave_readdata_5;
output 	rdclk_control_slave_readdata_6;
output 	rdclk_control_slave_readdata_7;
input 	wait_latency_counter_0;
input 	wait_latency_counter_1;
output 	wrfull;
output 	wrfull1;
output 	wrfull2;
input 	m0_write;
input 	in_data_reg_0;
input 	in_data_reg_1;
input 	in_data_reg_2;
input 	in_data_reg_3;
input 	in_data_reg_4;
input 	in_data_reg_5;
input 	in_data_reg_6;
input 	in_data_reg_7;
input 	in_data_reg_8;
input 	in_data_reg_9;
input 	in_data_reg_10;
input 	in_data_reg_11;
input 	in_data_reg_12;
input 	in_data_reg_13;
input 	in_data_reg_14;
input 	in_data_reg_15;
input 	in_data_reg_16;
input 	in_data_reg_17;
input 	in_data_reg_18;
input 	in_data_reg_19;
input 	in_data_reg_20;
input 	in_data_reg_21;
input 	in_data_reg_22;
input 	in_data_reg_23;
input 	in_data_reg_24;
input 	in_data_reg_25;
input 	in_data_reg_26;
input 	in_data_reg_27;
input 	in_data_reg_28;
input 	in_data_reg_29;
input 	in_data_reg_30;
input 	in_data_reg_31;
input 	r_sync_rst;
input 	r_sync_rst1;
input 	m0_write1;
input 	m0_read;
output 	wrclk_control_slave_readdata_0;
output 	wrclk_control_slave_readdata_1;
output 	wrclk_control_slave_readdata_2;
output 	wrclk_control_slave_readdata_3;
output 	wrclk_control_slave_readdata_4;
output 	wrclk_control_slave_readdata_5;
output 	wrclk_control_slave_readdata_6;
output 	wrclk_control_slave_readdata_7;
output 	wrfull3;
output 	wrfull4;
input 	int_nxt_addr_reg_dly_2;
input 	int_nxt_addr_reg_dly_4;
input 	int_nxt_addr_reg_dly_3;
input 	[31:0] wrclk_control_slave_writedata;
input 	in_data_reg_141;
input 	in_data_reg_81;
input 	in_data_reg_131;
input 	in_data_reg_121;
input 	in_data_reg_111;
input 	in_data_reg_101;
input 	in_data_reg_91;
input 	in_data_reg_191;
input 	in_data_reg_181;
input 	in_data_reg_171;
input 	in_data_reg_161;
input 	in_data_reg_151;
input 	in_data_reg_261;
input 	in_data_reg_211;
input 	in_data_reg_201;
input 	in_data_reg_311;
input 	in_data_reg_301;
input 	in_data_reg_291;
input 	in_data_reg_281;
input 	in_data_reg_271;
input 	in_data_reg_251;
input 	in_data_reg_241;
input 	in_data_reg_231;
input 	in_data_reg_221;
input 	in_data_reg_71;
input 	in_data_reg_61;
input 	fifo_hps_to_fpga_out_read;
input 	clock_bridge_0_in_clk_clk;
input 	fifo_hps_to_fpga_out_csr_address_2;
input 	fifo_hps_to_fpga_out_csr_address_0;
input 	fifo_hps_to_fpga_out_csr_address_1;
input 	fifo_hps_to_fpga_out_csr_read;
input 	[31:0] rdclk_control_slave_writedata;
input 	fifo_hps_to_fpga_out_csr_write;
input 	fifo_hps_to_fpga_out_csr_writedata_7;
input 	fifo_hps_to_fpga_out_csr_writedata_13;
input 	fifo_hps_to_fpga_out_csr_writedata_19;
input 	fifo_hps_to_fpga_out_csr_writedata_26;
input 	fifo_hps_to_fpga_out_csr_writedata_27;
input 	fifo_hps_to_fpga_out_csr_writedata_28;
input 	fifo_hps_to_fpga_out_csr_writedata_29;
input 	fifo_hps_to_fpga_out_csr_writedata_30;
input 	fifo_hps_to_fpga_out_csr_writedata_31;
input 	fifo_hps_to_fpga_out_csr_writedata_20;
input 	fifo_hps_to_fpga_out_csr_writedata_21;
input 	fifo_hps_to_fpga_out_csr_writedata_22;
input 	fifo_hps_to_fpga_out_csr_writedata_23;
input 	fifo_hps_to_fpga_out_csr_writedata_24;
input 	fifo_hps_to_fpga_out_csr_writedata_25;
input 	fifo_hps_to_fpga_out_csr_writedata_8;
input 	fifo_hps_to_fpga_out_csr_writedata_9;
input 	fifo_hps_to_fpga_out_csr_writedata_10;
input 	fifo_hps_to_fpga_out_csr_writedata_11;
input 	fifo_hps_to_fpga_out_csr_writedata_12;
input 	fifo_hps_to_fpga_out_csr_writedata_14;
input 	fifo_hps_to_fpga_out_csr_writedata_15;
input 	fifo_hps_to_fpga_out_csr_writedata_16;
input 	fifo_hps_to_fpga_out_csr_writedata_17;
input 	fifo_hps_to_fpga_out_csr_writedata_18;
input 	fifo_hps_to_fpga_out_csr_writedata_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_dcfifo|dual_clock_fifo|auto_generated|op_2~1_sumout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|op_2~5_sumout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|op_2~9_sumout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|op_2~17_sumout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|op_2~21_sumout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|op_1~1_sumout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|op_1~5_sumout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|op_1~9_sumout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|op_1~13_sumout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|op_1~17_sumout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|op_1~21_sumout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|op_1~25_sumout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|op_1~29_sumout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|rdempty_eq_comp|data_wire[2]~0_combout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|rdfull_eq_comp|aneb_result_wire[0]~0_combout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|rdfull_eq_comp|aneb_result_wire[0]~1_combout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~0_combout ;
wire \comb~0_combout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|rdfull_eq_comp|aneb_result_wire[0]~3_combout ;
wire \the_dcfifo|rdfull~0_combout ;
wire \the_dcfifo|rdfull~1_combout ;
wire \the_dcfifo|rdfull~2_combout ;
wire \wrdreq_sync_i|dreg[2]~q ;
wire \the_dcfifo|wrfull~7_combout ;
wire \the_dcfifo|dual_clock_fifo|auto_generated|wrempty_eq_comp|aneb_result_wire[0]~combout ;
wire \rdreq_sync_i|dreg[2]~q ;
wire \LessThan4~0_combout ;
wire \LessThan4~1_combout ;
wire \LessThan4~2_combout ;
wire \LessThan4~3_combout ;
wire \LessThan4~4_combout ;
wire \LessThan5~0_combout ;
wire \LessThan4~5_combout ;
wire \rdclk_control_slave_threshold_writedata[0]~0_combout ;
wire \rdclk_control_slave_almostempty_threshold_register[0]~0_combout ;
wire \always24~0_combout ;
wire \rdclk_control_slave_almostempty_threshold_register[0]~q ;
wire \rdclk_control_slave_status_full_q~q ;
wire \always32~0_combout ;
wire \rdclk_control_slave_full_n_reg~0_combout ;
wire \rdclk_control_slave_full_n_reg~q ;
wire \rdclk_control_slave_event_full_q~0_combout ;
wire \rdclk_control_slave_event_full_q~q ;
wire \always26~0_combout ;
wire \rdclk_control_slave_ienable_register[0]~q ;
wire \rdclk_control_slave_read_mux[0]~0_combout ;
wire \always25~0_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[0]~q ;
wire \rdclk_control_slave_read_mux[0]~28_combout ;
wire \rdclk_control_slave_threshold_writedata[1]~1_combout ;
wire \rdclk_control_slave_almostempty_threshold_register[1]~q ;
wire \rdclk_control_slave_status_empty_q~0_combout ;
wire \rdclk_control_slave_status_empty_q~q ;
wire \rdclk_control_slave_empty_n_reg~q ;
wire \rdclk_control_slave_event_empty_q~0_combout ;
wire \rdclk_control_slave_event_empty_q~1_combout ;
wire \rdclk_control_slave_event_empty_q~q ;
wire \rdclk_control_slave_ienable_register[1]~q ;
wire \rdclk_control_slave_read_mux[1]~1_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[1]~q ;
wire \rdclk_control_slave_read_mux[1]~24_combout ;
wire \LessThan5~1_combout ;
wire \rdclk_control_slave_threshold_writedata[2]~2_combout ;
wire \rdclk_control_slave_almostempty_threshold_register[2]~q ;
wire \rdclk_control_slave_threshold_writedata[6]~6_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[6]~4_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[6]~q ;
wire \rdclk_control_slave_threshold_writedata[7]~7_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[7]~5_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[7]~q ;
wire \rdclk_control_slave_threshold_writedata[5]~5_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[5]~3_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[5]~q ;
wire \LessThan7~0_combout ;
wire \rdclk_control_slave_threshold_writedata[4]~4_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[4]~2_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[4]~q ;
wire \LessThan7~1_combout ;
wire \rdclk_control_slave_threshold_writedata[3]~3_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[3]~1_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[3]~q ;
wire \LessThan7~2_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[2]~0_combout ;
wire \rdclk_control_slave_almostfull_threshold_register[2]~q ;
wire \LessThan7~3_combout ;
wire \LessThan7~4_combout ;
wire \LessThan7~5_combout ;
wire \LessThan7~6_combout ;
wire \rdclk_control_slave_status_almostfull_q~0_combout ;
wire \rdclk_control_slave_status_almostfull_q~q ;
wire \LessThan7~7_combout ;
wire \LessThan7~8_combout ;
wire \LessThan7~9_combout ;
wire \always30~0_combout ;
wire \rdclk_control_slave_almostfull_n_reg~q ;
wire \rdclk_control_slave_event_almostfull_q~0_combout ;
wire \rdclk_control_slave_event_almostfull_q~q ;
wire \rdclk_control_slave_ienable_register[2]~q ;
wire \rdclk_control_slave_read_mux[2]~2_combout ;
wire \rdclk_control_slave_read_mux[2]~20_combout ;
wire \rdclk_control_slave_almostempty_threshold_register[3]~q ;
wire \rdclk_control_slave_almostempty_threshold_register[6]~q ;
wire \rdclk_control_slave_almostempty_threshold_register[7]~q ;
wire \rdclk_control_slave_almostempty_threshold_register[5]~q ;
wire \LessThan6~0_combout ;
wire \rdclk_control_slave_almostempty_threshold_register[4]~q ;
wire \LessThan6~1_combout ;
wire \LessThan6~2_combout ;
wire \LessThan6~3_combout ;
wire \LessThan6~4_combout ;
wire \LessThan6~5_combout ;
wire \LessThan6~6_combout ;
wire \rdclk_control_slave_status_almostempty_q~0_combout ;
wire \rdclk_control_slave_status_almostempty_q~q ;
wire \LessThan6~7_combout ;
wire \LessThan6~8_combout ;
wire \LessThan6~9_combout ;
wire \always29~0_combout ;
wire \rdclk_control_slave_almostempty_n_reg~q ;
wire \rdclk_control_slave_event_almostempty_q~0_combout ;
wire \rdclk_control_slave_event_almostempty_q~q ;
wire \rdclk_control_slave_ienable_register[3]~q ;
wire \rdclk_control_slave_read_mux[3]~3_combout ;
wire \rdclk_control_slave_read_mux[3]~16_combout ;
wire \rdclk_control_slave_status_overflow_signal~combout ;
wire \rdclk_control_slave_status_overflow_q~q ;
wire \rdclk_control_slave_event_overflow_q~0_combout ;
wire \rdclk_control_slave_event_overflow_q~1_combout ;
wire \rdclk_control_slave_event_overflow_q~q ;
wire \rdclk_control_slave_ienable_register[4]~q ;
wire \rdclk_control_slave_read_mux[4]~4_combout ;
wire \rdclk_control_slave_read_mux[4]~12_combout ;
wire \rdclk_control_slave_status_underflow_signal~combout ;
wire \rdclk_control_slave_status_underflow_q~q ;
wire \always29~1_combout ;
wire \rdclk_control_slave_event_underflow_q~0_combout ;
wire \rdclk_control_slave_event_underflow_q~q ;
wire \rdclk_control_slave_ienable_register[5]~q ;
wire \rdclk_control_slave_read_mux[5]~5_combout ;
wire \rdclk_control_slave_read_mux[5]~8_combout ;
wire \rdclk_control_slave_read_mux[6]~6_combout ;
wire \rdclk_control_slave_read_mux[7]~7_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \LessThan0~2_combout ;
wire \LessThan0~3_combout ;
wire \LessThan0~4_combout ;
wire \LessThan0~5_combout ;
wire \LessThan1~0_combout ;
wire \wrclk_control_slave_threshold_writedata~0_combout ;
wire \LessThan0~6_combout ;
wire \LessThan0~7_combout ;
wire \wrclk_control_slave_threshold_writedata[0]~1_combout ;
wire \wrclk_control_slave_almostempty_threshold_register[0]~0_combout ;
wire \always4~0_combout ;
wire \always4~1_combout ;
wire \wrclk_control_slave_almostempty_threshold_register[0]~q ;
wire \wrclk_control_slave_status_full_q~q ;
wire \always7~0_combout ;
wire \wrclk_control_slave_full_n_reg~0_combout ;
wire \wrclk_control_slave_full_n_reg~q ;
wire \wrclk_control_slave_event_full_q~0_combout ;
wire \wrclk_control_slave_event_full_q~q ;
wire \always6~0_combout ;
wire \wrclk_control_slave_ienable_register[0]~q ;
wire \wrclk_control_slave_read_mux[0]~0_combout ;
wire \always5~0_combout ;
wire \wrclk_control_slave_almostfull_threshold_register[0]~q ;
wire \wrclk_control_slave_read_mux[0]~28_combout ;
wire \wrclk_control_slave_threshold_writedata[1]~2_combout ;
wire \wrclk_control_slave_almostempty_threshold_register[1]~q ;
wire \wrclk_control_slave_status_empty_q~0_combout ;
wire \wrclk_control_slave_status_empty_q~q ;
wire \wrclk_control_slave_empty_n_reg~q ;
wire \wrclk_control_slave_event_empty_q~0_combout ;
wire \wrclk_control_slave_event_empty_q~q ;
wire \wrclk_control_slave_ienable_register[1]~q ;
wire \wrclk_control_slave_read_mux[1]~1_combout ;
wire \wrclk_control_slave_almostfull_threshold_register[1]~q ;
wire \wrclk_control_slave_read_mux[1]~24_combout ;
wire \wrclk_control_slave_threshold_writedata[2]~3_combout ;
wire \wrclk_control_slave_almostempty_threshold_register[2]~q ;
wire \wrclk_control_slave_almostfull_threshold_register[2]~0_combout ;
wire \wrclk_control_slave_almostfull_threshold_register[2]~q ;
wire \wrclk_control_slave_threshold_writedata[3]~4_combout ;
wire \wrclk_control_slave_almostfull_threshold_register[3]~1_combout ;
wire \wrclk_control_slave_almostfull_threshold_register[3]~q ;
wire \LessThan3~0_combout ;
wire \LessThan3~2_combout ;
wire \wrclk_control_slave_threshold_writedata[6]~7_combout ;
wire \wrclk_control_slave_almostfull_threshold_register[6]~4_combout ;
wire \wrclk_control_slave_almostfull_threshold_register[6]~q ;
wire \wrclk_control_slave_threshold_writedata[4]~5_combout ;
wire \wrclk_control_slave_almostfull_threshold_register[4]~2_combout ;
wire \wrclk_control_slave_almostfull_threshold_register[4]~q ;
wire \LessThan3~3_combout ;
wire \wrclk_control_slave_threshold_writedata[7]~8_combout ;
wire \wrclk_control_slave_almostfull_threshold_register[7]~5_combout ;
wire \wrclk_control_slave_almostfull_threshold_register[7]~q ;
wire \wrclk_control_slave_threshold_writedata[5]~6_combout ;
wire \wrclk_control_slave_almostfull_threshold_register[5]~3_combout ;
wire \wrclk_control_slave_almostfull_threshold_register[5]~q ;
wire \LessThan3~4_combout ;
wire \LessThan3~5_combout ;
wire \LessThan3~1_combout ;
wire \wrclk_control_slave_status_almostfull_q~0_combout ;
wire \wrclk_control_slave_status_almostfull_q~q ;
wire \wrclk_control_slave_almostfull_n_reg~q ;
wire \wrclk_control_slave_event_almostfull_q~0_combout ;
wire \wrclk_control_slave_event_almostfull_q~q ;
wire \wrclk_control_slave_ienable_register[2]~q ;
wire \wrclk_control_slave_read_mux[2]~2_combout ;
wire \wrclk_control_slave_read_mux[2]~20_combout ;
wire \wrclk_control_slave_almostempty_threshold_register[3]~q ;
wire \LessThan2~0_combout ;
wire \LessThan2~2_combout ;
wire \wrclk_control_slave_almostempty_threshold_register[6]~q ;
wire \wrclk_control_slave_almostempty_threshold_register[4]~q ;
wire \LessThan2~3_combout ;
wire \wrclk_control_slave_almostempty_threshold_register[7]~q ;
wire \wrclk_control_slave_almostempty_threshold_register[5]~q ;
wire \LessThan2~4_combout ;
wire \LessThan2~5_combout ;
wire \LessThan2~1_combout ;
wire \wrclk_control_slave_status_almostempty_q~0_combout ;
wire \wrclk_control_slave_status_almostempty_q~q ;
wire \wrclk_control_slave_almostempty_n_reg~q ;
wire \wrclk_control_slave_event_almostempty_q~0_combout ;
wire \wrclk_control_slave_event_almostempty_q~q ;
wire \wrclk_control_slave_ienable_register[3]~q ;
wire \wrclk_control_slave_read_mux[3]~3_combout ;
wire \wrclk_control_slave_read_mux[3]~16_combout ;
wire \wrclk_control_slave_status_overflow_signal~combout ;
wire \wrclk_control_slave_status_overflow_q~q ;
wire \wrclk_control_slave_event_overflow_q~0_combout ;
wire \wrclk_control_slave_event_overflow_q~q ;
wire \wrclk_control_slave_ienable_register[4]~q ;
wire \wrclk_control_slave_read_mux[4]~4_combout ;
wire \wrclk_control_slave_read_mux[4]~12_combout ;
wire \wrclk_control_slave_status_underflow_signal~combout ;
wire \wrclk_control_slave_status_underflow_q~q ;
wire \wrclk_control_slave_event_underflow_q~0_combout ;
wire \wrclk_control_slave_event_underflow_q~q ;
wire \wrclk_control_slave_ienable_register[5]~q ;
wire \wrclk_control_slave_read_mux[5]~5_combout ;
wire \wrclk_control_slave_read_mux[5]~8_combout ;
wire \wrclk_control_slave_read_mux[6]~6_combout ;
wire \wrclk_control_slave_read_mux[7]~7_combout ;


Computer_System_altera_std_synchronizer_1 wrdreq_sync_i(
	.din(m0_write),
	.reset_n(r_sync_rst),
	.dreg_2(\wrdreq_sync_i|dreg[2]~q ),
	.clk(clock_bridge_0_in_clk_clk));

Computer_System_altera_std_synchronizer rdreq_sync_i(
	.clk(outclk_wire_0),
	.reset_n(r_sync_rst1),
	.dreg_2(\rdreq_sync_i|dreg[2]~q ),
	.din(fifo_hps_to_fpga_out_read));

Computer_System_Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo the_dcfifo(
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.outclk_wire_0(outclk_wire_0),
	.op_2(\the_dcfifo|dual_clock_fifo|auto_generated|op_2~1_sumout ),
	.op_21(\the_dcfifo|dual_clock_fifo|auto_generated|op_2~5_sumout ),
	.op_22(\the_dcfifo|dual_clock_fifo|auto_generated|op_2~9_sumout ),
	.op_23(op_2),
	.op_24(\the_dcfifo|dual_clock_fifo|auto_generated|op_2~17_sumout ),
	.op_25(\the_dcfifo|dual_clock_fifo|auto_generated|op_2~21_sumout ),
	.op_26(op_21),
	.op_27(op_22),
	.op_1(\the_dcfifo|dual_clock_fifo|auto_generated|op_1~1_sumout ),
	.op_11(\the_dcfifo|dual_clock_fifo|auto_generated|op_1~5_sumout ),
	.op_12(\the_dcfifo|dual_clock_fifo|auto_generated|op_1~9_sumout ),
	.op_13(\the_dcfifo|dual_clock_fifo|auto_generated|op_1~13_sumout ),
	.op_14(\the_dcfifo|dual_clock_fifo|auto_generated|op_1~17_sumout ),
	.op_15(\the_dcfifo|dual_clock_fifo|auto_generated|op_1~21_sumout ),
	.op_16(\the_dcfifo|dual_clock_fifo|auto_generated|op_1~25_sumout ),
	.op_17(\the_dcfifo|dual_clock_fifo|auto_generated|op_1~29_sumout ),
	.data_wire_2(\the_dcfifo|dual_clock_fifo|auto_generated|rdempty_eq_comp|data_wire[2]~0_combout ),
	.aneb_result_wire_0(\the_dcfifo|dual_clock_fifo|auto_generated|rdfull_eq_comp|aneb_result_wire[0]~0_combout ),
	.aneb_result_wire_01(\the_dcfifo|dual_clock_fifo|auto_generated|rdfull_eq_comp|aneb_result_wire[0]~1_combout ),
	.aneb_result_wire_02(\the_dcfifo|dual_clock_fifo|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~0_combout ),
	.aneb_result_wire_03(aneb_result_wire_0),
	.wrfull(wrfull),
	.wrfull1(wrfull1),
	.wrfull2(wrfull2),
	.m0_write(m0_write),
	.in_data_reg_0(in_data_reg_0),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_24(in_data_reg_24),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_31(in_data_reg_31),
	.wrfull3(wrfull3),
	.wrfull4(wrfull4),
	.comb(\comb~0_combout ),
	.aneb_result_wire_04(\the_dcfifo|dual_clock_fifo|auto_generated|rdfull_eq_comp|aneb_result_wire[0]~3_combout ),
	.rdfull(\the_dcfifo|rdfull~0_combout ),
	.rdfull1(\the_dcfifo|rdfull~1_combout ),
	.rdfull2(\the_dcfifo|rdfull~2_combout ),
	.wrfull5(\the_dcfifo|wrfull~7_combout ),
	.aneb_result_wire_05(\the_dcfifo|dual_clock_fifo|auto_generated|wrempty_eq_comp|aneb_result_wire[0]~combout ),
	.fifo_hps_to_fpga_out_read(fifo_hps_to_fpga_out_read),
	.clock_bridge_0_in_clk_clk(clock_bridge_0_in_clk_clk));

cyclonev_lcell_comb \comb~0 (
	.dataa(!r_sync_rst),
	.datab(!r_sync_rst1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h7777777777777777;
defparam \comb~0 .shared_arith = "off";

dffeas \rdclk_control_slave_readdata[0] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_read_mux[0]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_hps_to_fpga_out_csr_read),
	.q(rdclk_control_slave_readdata_0),
	.prn(vcc));
defparam \rdclk_control_slave_readdata[0] .is_wysiwyg = "true";
defparam \rdclk_control_slave_readdata[0] .power_up = "low";

dffeas \rdclk_control_slave_readdata[1] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_read_mux[1]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_hps_to_fpga_out_csr_read),
	.q(rdclk_control_slave_readdata_1),
	.prn(vcc));
defparam \rdclk_control_slave_readdata[1] .is_wysiwyg = "true";
defparam \rdclk_control_slave_readdata[1] .power_up = "low";

dffeas \rdclk_control_slave_readdata[2] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_read_mux[2]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_hps_to_fpga_out_csr_read),
	.q(rdclk_control_slave_readdata_2),
	.prn(vcc));
defparam \rdclk_control_slave_readdata[2] .is_wysiwyg = "true";
defparam \rdclk_control_slave_readdata[2] .power_up = "low";

dffeas \rdclk_control_slave_readdata[3] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_read_mux[3]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_hps_to_fpga_out_csr_read),
	.q(rdclk_control_slave_readdata_3),
	.prn(vcc));
defparam \rdclk_control_slave_readdata[3] .is_wysiwyg = "true";
defparam \rdclk_control_slave_readdata[3] .power_up = "low";

dffeas \rdclk_control_slave_readdata[4] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_read_mux[4]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_hps_to_fpga_out_csr_read),
	.q(rdclk_control_slave_readdata_4),
	.prn(vcc));
defparam \rdclk_control_slave_readdata[4] .is_wysiwyg = "true";
defparam \rdclk_control_slave_readdata[4] .power_up = "low";

dffeas \rdclk_control_slave_readdata[5] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_read_mux[5]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_hps_to_fpga_out_csr_read),
	.q(rdclk_control_slave_readdata_5),
	.prn(vcc));
defparam \rdclk_control_slave_readdata[5] .is_wysiwyg = "true";
defparam \rdclk_control_slave_readdata[5] .power_up = "low";

dffeas \rdclk_control_slave_readdata[6] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_read_mux[6]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_hps_to_fpga_out_csr_read),
	.q(rdclk_control_slave_readdata_6),
	.prn(vcc));
defparam \rdclk_control_slave_readdata[6] .is_wysiwyg = "true";
defparam \rdclk_control_slave_readdata[6] .power_up = "low";

dffeas \rdclk_control_slave_readdata[7] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_read_mux[7]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_hps_to_fpga_out_csr_read),
	.q(rdclk_control_slave_readdata_7),
	.prn(vcc));
defparam \rdclk_control_slave_readdata[7] .is_wysiwyg = "true";
defparam \rdclk_control_slave_readdata[7] .power_up = "low";

dffeas \wrclk_control_slave_readdata[0] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_read_mux[0]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(m0_read),
	.q(wrclk_control_slave_readdata_0),
	.prn(vcc));
defparam \wrclk_control_slave_readdata[0] .is_wysiwyg = "true";
defparam \wrclk_control_slave_readdata[0] .power_up = "low";

dffeas \wrclk_control_slave_readdata[1] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_read_mux[1]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(m0_read),
	.q(wrclk_control_slave_readdata_1),
	.prn(vcc));
defparam \wrclk_control_slave_readdata[1] .is_wysiwyg = "true";
defparam \wrclk_control_slave_readdata[1] .power_up = "low";

dffeas \wrclk_control_slave_readdata[2] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_read_mux[2]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(m0_read),
	.q(wrclk_control_slave_readdata_2),
	.prn(vcc));
defparam \wrclk_control_slave_readdata[2] .is_wysiwyg = "true";
defparam \wrclk_control_slave_readdata[2] .power_up = "low";

dffeas \wrclk_control_slave_readdata[3] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_read_mux[3]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(m0_read),
	.q(wrclk_control_slave_readdata_3),
	.prn(vcc));
defparam \wrclk_control_slave_readdata[3] .is_wysiwyg = "true";
defparam \wrclk_control_slave_readdata[3] .power_up = "low";

dffeas \wrclk_control_slave_readdata[4] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_read_mux[4]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(m0_read),
	.q(wrclk_control_slave_readdata_4),
	.prn(vcc));
defparam \wrclk_control_slave_readdata[4] .is_wysiwyg = "true";
defparam \wrclk_control_slave_readdata[4] .power_up = "low";

dffeas \wrclk_control_slave_readdata[5] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_read_mux[5]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(m0_read),
	.q(wrclk_control_slave_readdata_5),
	.prn(vcc));
defparam \wrclk_control_slave_readdata[5] .is_wysiwyg = "true";
defparam \wrclk_control_slave_readdata[5] .power_up = "low";

dffeas \wrclk_control_slave_readdata[6] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_read_mux[6]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(m0_read),
	.q(wrclk_control_slave_readdata_6),
	.prn(vcc));
defparam \wrclk_control_slave_readdata[6] .is_wysiwyg = "true";
defparam \wrclk_control_slave_readdata[6] .power_up = "low";

dffeas \wrclk_control_slave_readdata[7] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_read_mux[7]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(m0_read),
	.q(wrclk_control_slave_readdata_7),
	.prn(vcc));
defparam \wrclk_control_slave_readdata[7] .is_wysiwyg = "true";
defparam \wrclk_control_slave_readdata[7] .power_up = "low";

cyclonev_lcell_comb \LessThan4~0 (
	.dataa(!fifo_hps_to_fpga_out_csr_writedata_26),
	.datab(!fifo_hps_to_fpga_out_csr_writedata_27),
	.datac(!fifo_hps_to_fpga_out_csr_writedata_28),
	.datad(!fifo_hps_to_fpga_out_csr_writedata_29),
	.datae(!fifo_hps_to_fpga_out_csr_writedata_30),
	.dataf(!fifo_hps_to_fpga_out_csr_writedata_31),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~0 .extended_lut = "off";
defparam \LessThan4~0 .lut_mask = 64'h8000000000000000;
defparam \LessThan4~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~1 (
	.dataa(!fifo_hps_to_fpga_out_csr_writedata_20),
	.datab(!fifo_hps_to_fpga_out_csr_writedata_21),
	.datac(!fifo_hps_to_fpga_out_csr_writedata_22),
	.datad(!fifo_hps_to_fpga_out_csr_writedata_23),
	.datae(!fifo_hps_to_fpga_out_csr_writedata_24),
	.dataf(!fifo_hps_to_fpga_out_csr_writedata_25),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~1 .extended_lut = "off";
defparam \LessThan4~1 .lut_mask = 64'h8000000000000000;
defparam \LessThan4~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~2 (
	.dataa(!fifo_hps_to_fpga_out_csr_writedata_8),
	.datab(!fifo_hps_to_fpga_out_csr_writedata_9),
	.datac(!fifo_hps_to_fpga_out_csr_writedata_10),
	.datad(!fifo_hps_to_fpga_out_csr_writedata_11),
	.datae(!fifo_hps_to_fpga_out_csr_writedata_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~2 .extended_lut = "off";
defparam \LessThan4~2 .lut_mask = 64'h8000000080000000;
defparam \LessThan4~2 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~3 (
	.dataa(!fifo_hps_to_fpga_out_csr_writedata_14),
	.datab(!fifo_hps_to_fpga_out_csr_writedata_15),
	.datac(!fifo_hps_to_fpga_out_csr_writedata_16),
	.datad(!fifo_hps_to_fpga_out_csr_writedata_17),
	.datae(!fifo_hps_to_fpga_out_csr_writedata_18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~3 .extended_lut = "off";
defparam \LessThan4~3 .lut_mask = 64'h8000000080000000;
defparam \LessThan4~3 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~4 (
	.dataa(!fifo_hps_to_fpga_out_csr_writedata_13),
	.datab(!fifo_hps_to_fpga_out_csr_writedata_19),
	.datac(!\LessThan4~0_combout ),
	.datad(!\LessThan4~1_combout ),
	.datae(!\LessThan4~2_combout ),
	.dataf(!\LessThan4~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~4 .extended_lut = "off";
defparam \LessThan4~4 .lut_mask = 64'h0000000000000008;
defparam \LessThan4~4 .shared_arith = "off";

cyclonev_lcell_comb \LessThan5~0 (
	.dataa(!rdclk_control_slave_writedata[2]),
	.datab(!rdclk_control_slave_writedata[3]),
	.datac(!rdclk_control_slave_writedata[4]),
	.datad(!rdclk_control_slave_writedata[5]),
	.datae(!fifo_hps_to_fpga_out_csr_writedata_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan5~0 .extended_lut = "off";
defparam \LessThan5~0 .lut_mask = 64'h0000000100000001;
defparam \LessThan5~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~5 (
	.dataa(!rdclk_control_slave_writedata[2]),
	.datab(!rdclk_control_slave_writedata[3]),
	.datac(!rdclk_control_slave_writedata[4]),
	.datad(!rdclk_control_slave_writedata[5]),
	.datae(!fifo_hps_to_fpga_out_csr_writedata_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~5 .extended_lut = "off";
defparam \LessThan4~5 .lut_mask = 64'h8000000080000000;
defparam \LessThan4~5 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_threshold_writedata[0]~0 (
	.dataa(!rdclk_control_slave_writedata[0]),
	.datab(!fifo_hps_to_fpga_out_csr_writedata_7),
	.datac(!rdclk_control_slave_writedata[1]),
	.datad(!\LessThan4~4_combout ),
	.datae(!\LessThan5~0_combout ),
	.dataf(!\LessThan4~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_threshold_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_threshold_writedata[0]~0 .extended_lut = "off";
defparam \rdclk_control_slave_threshold_writedata[0]~0 .lut_mask = 64'h0055004400D500C4;
defparam \rdclk_control_slave_threshold_writedata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_almostempty_threshold_register[0]~0 (
	.dataa(!\rdclk_control_slave_threshold_writedata[0]~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_almostempty_threshold_register[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_almostempty_threshold_register[0]~0 .extended_lut = "off";
defparam \rdclk_control_slave_almostempty_threshold_register[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdclk_control_slave_almostempty_threshold_register[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \always24~0 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!fifo_hps_to_fpga_out_csr_write),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always24~0 .extended_lut = "off";
defparam \always24~0 .lut_mask = 64'h0010001000100010;
defparam \always24~0 .shared_arith = "off";

dffeas \rdclk_control_slave_almostempty_threshold_register[0] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_almostempty_threshold_register[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always24~0_combout ),
	.q(\rdclk_control_slave_almostempty_threshold_register[0]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostempty_threshold_register[0] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostempty_threshold_register[0] .power_up = "low";

dffeas rdclk_control_slave_status_full_q(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\the_dcfifo|rdfull~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_status_full_q~q ),
	.prn(vcc));
defparam rdclk_control_slave_status_full_q.is_wysiwyg = "true";
defparam rdclk_control_slave_status_full_q.power_up = "low";

cyclonev_lcell_comb \always32~0 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!rdclk_control_slave_writedata[0]),
	.datae(!fifo_hps_to_fpga_out_csr_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always32~0 .extended_lut = "off";
defparam \always32~0 .lut_mask = 64'h0000000800000008;
defparam \always32~0 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_full_n_reg~0 (
	.dataa(!\the_dcfifo|rdfull~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_full_n_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_full_n_reg~0 .extended_lut = "off";
defparam \rdclk_control_slave_full_n_reg~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdclk_control_slave_full_n_reg~0 .shared_arith = "off";

dffeas rdclk_control_slave_full_n_reg(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_full_n_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_full_n_reg~q ),
	.prn(vcc));
defparam rdclk_control_slave_full_n_reg.is_wysiwyg = "true";
defparam rdclk_control_slave_full_n_reg.power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_event_full_q~0 (
	.dataa(!\rdclk_control_slave_event_full_q~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|rdfull_eq_comp|aneb_result_wire[0]~3_combout ),
	.datac(!\the_dcfifo|rdfull~0_combout ),
	.datad(!\the_dcfifo|rdfull~1_combout ),
	.datae(!\always32~0_combout ),
	.dataf(!\rdclk_control_slave_full_n_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_event_full_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_event_full_q~0 .extended_lut = "off";
defparam \rdclk_control_slave_event_full_q~0 .lut_mask = 64'h55550000777F0000;
defparam \rdclk_control_slave_event_full_q~0 .shared_arith = "off";

dffeas rdclk_control_slave_event_full_q(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_event_full_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_event_full_q~q ),
	.prn(vcc));
defparam rdclk_control_slave_event_full_q.is_wysiwyg = "true";
defparam rdclk_control_slave_event_full_q.power_up = "low";

cyclonev_lcell_comb \always26~0 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!fifo_hps_to_fpga_out_csr_write),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always26~0 .extended_lut = "off";
defparam \always26~0 .lut_mask = 64'h0002000200020002;
defparam \always26~0 .shared_arith = "off";

dffeas \rdclk_control_slave_ienable_register[0] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(rdclk_control_slave_writedata[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always26~0_combout ),
	.q(\rdclk_control_slave_ienable_register[0]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_ienable_register[0] .is_wysiwyg = "true";
defparam \rdclk_control_slave_ienable_register[0] .power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[0]~0 (
	.dataa(!\rdclk_control_slave_status_full_q~q ),
	.datab(!fifo_hps_to_fpga_out_csr_address_2),
	.datac(!fifo_hps_to_fpga_out_csr_address_0),
	.datad(!fifo_hps_to_fpga_out_csr_address_1),
	.datae(!\rdclk_control_slave_event_full_q~q ),
	.dataf(!\rdclk_control_slave_ienable_register[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[0]~0 .extended_lut = "off";
defparam \rdclk_control_slave_read_mux[0]~0 .lut_mask = 64'h040004C0040C04CC;
defparam \rdclk_control_slave_read_mux[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \always25~0 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!fifo_hps_to_fpga_out_csr_write),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always25~0 .extended_lut = "off";
defparam \always25~0 .lut_mask = 64'h0040004000400040;
defparam \always25~0 .shared_arith = "off";

dffeas \rdclk_control_slave_almostfull_threshold_register[0] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_threshold_writedata[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always25~0_combout ),
	.q(\rdclk_control_slave_almostfull_threshold_register[0]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostfull_threshold_register[0] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostfull_threshold_register[0] .power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[0]~28 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_1),
	.datab(!fifo_hps_to_fpga_out_csr_address_2),
	.datac(!\rdclk_control_slave_almostempty_threshold_register[0]~q ),
	.datad(!\rdclk_control_slave_read_mux[0]~0_combout ),
	.datae(!fifo_hps_to_fpga_out_csr_address_0),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~1_sumout ),
	.datag(!\rdclk_control_slave_almostfull_threshold_register[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[0]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[0]~28 .extended_lut = "on";
defparam \rdclk_control_slave_read_mux[0]~28 .lut_mask = 64'h02FF20FF9BFF31FF;
defparam \rdclk_control_slave_read_mux[0]~28 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_threshold_writedata[1]~1 (
	.dataa(gnd),
	.datab(!fifo_hps_to_fpga_out_csr_writedata_7),
	.datac(!rdclk_control_slave_writedata[1]),
	.datad(!\LessThan4~4_combout ),
	.datae(!\LessThan5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_threshold_writedata[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_threshold_writedata[1]~1 .extended_lut = "off";
defparam \rdclk_control_slave_threshold_writedata[1]~1 .lut_mask = 64'h000F000C000F000C;
defparam \rdclk_control_slave_threshold_writedata[1]~1 .shared_arith = "off";

dffeas \rdclk_control_slave_almostempty_threshold_register[1] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_threshold_writedata[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always24~0_combout ),
	.q(\rdclk_control_slave_almostempty_threshold_register[1]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostempty_threshold_register[1] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostempty_threshold_register[1] .power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_status_empty_q~0 (
	.dataa(!aneb_result_wire_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_status_empty_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_status_empty_q~0 .extended_lut = "off";
defparam \rdclk_control_slave_status_empty_q~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdclk_control_slave_status_empty_q~0 .shared_arith = "off";

dffeas rdclk_control_slave_status_empty_q(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_status_empty_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_status_empty_q~q ),
	.prn(vcc));
defparam rdclk_control_slave_status_empty_q.is_wysiwyg = "true";
defparam rdclk_control_slave_status_empty_q.power_up = "low";

dffeas rdclk_control_slave_empty_n_reg(
	.clk(clock_bridge_0_in_clk_clk),
	.d(aneb_result_wire_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_empty_n_reg~q ),
	.prn(vcc));
defparam rdclk_control_slave_empty_n_reg.is_wysiwyg = "true";
defparam rdclk_control_slave_empty_n_reg.power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_event_empty_q~0 (
	.dataa(!\the_dcfifo|dual_clock_fifo|auto_generated|rdempty_eq_comp|data_wire[2]~0_combout ),
	.datab(!\rdclk_control_slave_event_empty_q~q ),
	.datac(!\the_dcfifo|dual_clock_fifo|auto_generated|rdfull_eq_comp|aneb_result_wire[0]~0_combout ),
	.datad(!\the_dcfifo|dual_clock_fifo|auto_generated|rdfull_eq_comp|aneb_result_wire[0]~1_combout ),
	.datae(!\the_dcfifo|dual_clock_fifo|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~0_combout ),
	.dataf(!\rdclk_control_slave_empty_n_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_event_empty_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_event_empty_q~0 .extended_lut = "off";
defparam \rdclk_control_slave_event_empty_q~0 .lut_mask = 64'hCCCCCCCCCCCCCCC4;
defparam \rdclk_control_slave_event_empty_q~0 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_event_empty_q~1 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!fifo_hps_to_fpga_out_csr_write),
	.datae(!rdclk_control_slave_writedata[1]),
	.dataf(!\rdclk_control_slave_event_empty_q~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_event_empty_q~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_event_empty_q~1 .extended_lut = "off";
defparam \rdclk_control_slave_event_empty_q~1 .lut_mask = 64'hFFFFFFF700000000;
defparam \rdclk_control_slave_event_empty_q~1 .shared_arith = "off";

dffeas rdclk_control_slave_event_empty_q(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_event_empty_q~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_event_empty_q~q ),
	.prn(vcc));
defparam rdclk_control_slave_event_empty_q.is_wysiwyg = "true";
defparam rdclk_control_slave_event_empty_q.power_up = "low";

dffeas \rdclk_control_slave_ienable_register[1] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(rdclk_control_slave_writedata[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always26~0_combout ),
	.q(\rdclk_control_slave_ienable_register[1]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_ienable_register[1] .is_wysiwyg = "true";
defparam \rdclk_control_slave_ienable_register[1] .power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[1]~1 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!\rdclk_control_slave_status_empty_q~q ),
	.datae(!\rdclk_control_slave_event_empty_q~q ),
	.dataf(!\rdclk_control_slave_ienable_register[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[1]~1 .extended_lut = "off";
defparam \rdclk_control_slave_read_mux[1]~1 .lut_mask = 64'h0020082802220A2A;
defparam \rdclk_control_slave_read_mux[1]~1 .shared_arith = "off";

dffeas \rdclk_control_slave_almostfull_threshold_register[1] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_threshold_writedata[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always25~0_combout ),
	.q(\rdclk_control_slave_almostfull_threshold_register[1]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostfull_threshold_register[1] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostfull_threshold_register[1] .power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[1]~24 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_1),
	.datab(!fifo_hps_to_fpga_out_csr_address_2),
	.datac(!\rdclk_control_slave_almostempty_threshold_register[1]~q ),
	.datad(!\rdclk_control_slave_read_mux[1]~1_combout ),
	.datae(!fifo_hps_to_fpga_out_csr_address_0),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~5_sumout ),
	.datag(!\rdclk_control_slave_almostfull_threshold_register[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[1]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[1]~24 .extended_lut = "on";
defparam \rdclk_control_slave_read_mux[1]~24 .lut_mask = 64'h02FF02FF9BFF13FF;
defparam \rdclk_control_slave_read_mux[1]~24 .shared_arith = "off";

cyclonev_lcell_comb \LessThan5~1 (
	.dataa(!rdclk_control_slave_writedata[0]),
	.datab(!rdclk_control_slave_writedata[1]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan5~1 .extended_lut = "off";
defparam \LessThan5~1 .lut_mask = 64'h8888888888888888;
defparam \LessThan5~1 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_threshold_writedata[2]~2 (
	.dataa(!rdclk_control_slave_writedata[2]),
	.datab(!fifo_hps_to_fpga_out_csr_writedata_7),
	.datac(!\LessThan5~1_combout ),
	.datad(!\LessThan4~4_combout ),
	.datae(!\LessThan5~0_combout ),
	.dataf(!\LessThan4~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_threshold_writedata[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_threshold_writedata[2]~2 .extended_lut = "off";
defparam \rdclk_control_slave_threshold_writedata[2]~2 .lut_mask = 64'hFF55FF75FF51FF71;
defparam \rdclk_control_slave_threshold_writedata[2]~2 .shared_arith = "off";

dffeas \rdclk_control_slave_almostempty_threshold_register[2] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_threshold_writedata[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always24~0_combout ),
	.q(\rdclk_control_slave_almostempty_threshold_register[2]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostempty_threshold_register[2] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostempty_threshold_register[2] .power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_threshold_writedata[6]~6 (
	.dataa(!fifo_hps_to_fpga_out_csr_writedata_6),
	.datab(!fifo_hps_to_fpga_out_csr_writedata_7),
	.datac(!\LessThan5~1_combout ),
	.datad(!\LessThan4~4_combout ),
	.datae(!\LessThan5~0_combout ),
	.dataf(!\LessThan4~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_threshold_writedata[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_threshold_writedata[6]~6 .extended_lut = "off";
defparam \rdclk_control_slave_threshold_writedata[6]~6 .lut_mask = 64'hFF55FF75FF51FF71;
defparam \rdclk_control_slave_threshold_writedata[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_almostfull_threshold_register[6]~4 (
	.dataa(!\rdclk_control_slave_threshold_writedata[6]~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_almostfull_threshold_register[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_almostfull_threshold_register[6]~4 .extended_lut = "off";
defparam \rdclk_control_slave_almostfull_threshold_register[6]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdclk_control_slave_almostfull_threshold_register[6]~4 .shared_arith = "off";

dffeas \rdclk_control_slave_almostfull_threshold_register[6] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_almostfull_threshold_register[6]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always25~0_combout ),
	.q(\rdclk_control_slave_almostfull_threshold_register[6]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostfull_threshold_register[6] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostfull_threshold_register[6] .power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_threshold_writedata[7]~7 (
	.dataa(!fifo_hps_to_fpga_out_csr_writedata_7),
	.datab(gnd),
	.datac(!\LessThan4~4_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_threshold_writedata[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_threshold_writedata[7]~7 .extended_lut = "off";
defparam \rdclk_control_slave_threshold_writedata[7]~7 .lut_mask = 64'hF5F5F5F5F5F5F5F5;
defparam \rdclk_control_slave_threshold_writedata[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_almostfull_threshold_register[7]~5 (
	.dataa(!\rdclk_control_slave_threshold_writedata[7]~7_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_almostfull_threshold_register[7]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_almostfull_threshold_register[7]~5 .extended_lut = "off";
defparam \rdclk_control_slave_almostfull_threshold_register[7]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdclk_control_slave_almostfull_threshold_register[7]~5 .shared_arith = "off";

dffeas \rdclk_control_slave_almostfull_threshold_register[7] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_almostfull_threshold_register[7]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always25~0_combout ),
	.q(\rdclk_control_slave_almostfull_threshold_register[7]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostfull_threshold_register[7] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostfull_threshold_register[7] .power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_threshold_writedata[5]~5 (
	.dataa(!rdclk_control_slave_writedata[5]),
	.datab(!fifo_hps_to_fpga_out_csr_writedata_7),
	.datac(!\LessThan5~1_combout ),
	.datad(!\LessThan4~4_combout ),
	.datae(!\LessThan5~0_combout ),
	.dataf(!\LessThan4~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_threshold_writedata[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_threshold_writedata[5]~5 .extended_lut = "off";
defparam \rdclk_control_slave_threshold_writedata[5]~5 .lut_mask = 64'hFF55FF75FF51FF71;
defparam \rdclk_control_slave_threshold_writedata[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_almostfull_threshold_register[5]~3 (
	.dataa(!\rdclk_control_slave_threshold_writedata[5]~5_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_almostfull_threshold_register[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_almostfull_threshold_register[5]~3 .extended_lut = "off";
defparam \rdclk_control_slave_almostfull_threshold_register[5]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdclk_control_slave_almostfull_threshold_register[5]~3 .shared_arith = "off";

dffeas \rdclk_control_slave_almostfull_threshold_register[5] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_almostfull_threshold_register[5]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always25~0_combout ),
	.q(\rdclk_control_slave_almostfull_threshold_register[5]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostfull_threshold_register[5] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostfull_threshold_register[5] .power_up = "low";

cyclonev_lcell_comb \LessThan7~0 (
	.dataa(!\rdclk_control_slave_almostfull_threshold_register[5]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~21_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan7~0 .extended_lut = "off";
defparam \LessThan7~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan7~0 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_threshold_writedata[4]~4 (
	.dataa(!rdclk_control_slave_writedata[4]),
	.datab(!fifo_hps_to_fpga_out_csr_writedata_7),
	.datac(!\LessThan5~1_combout ),
	.datad(!\LessThan4~4_combout ),
	.datae(!\LessThan5~0_combout ),
	.dataf(!\LessThan4~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_threshold_writedata[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_threshold_writedata[4]~4 .extended_lut = "off";
defparam \rdclk_control_slave_threshold_writedata[4]~4 .lut_mask = 64'hFF55FF75FF51FF71;
defparam \rdclk_control_slave_threshold_writedata[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_almostfull_threshold_register[4]~2 (
	.dataa(!\rdclk_control_slave_threshold_writedata[4]~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_almostfull_threshold_register[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_almostfull_threshold_register[4]~2 .extended_lut = "off";
defparam \rdclk_control_slave_almostfull_threshold_register[4]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdclk_control_slave_almostfull_threshold_register[4]~2 .shared_arith = "off";

dffeas \rdclk_control_slave_almostfull_threshold_register[4] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_almostfull_threshold_register[4]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always25~0_combout ),
	.q(\rdclk_control_slave_almostfull_threshold_register[4]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostfull_threshold_register[4] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostfull_threshold_register[4] .power_up = "low";

cyclonev_lcell_comb \LessThan7~1 (
	.dataa(!\rdclk_control_slave_almostfull_threshold_register[5]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~21_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan7~1 .extended_lut = "off";
defparam \LessThan7~1 .lut_mask = 64'h6666666666666666;
defparam \LessThan7~1 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_threshold_writedata[3]~3 (
	.dataa(!rdclk_control_slave_writedata[3]),
	.datab(!fifo_hps_to_fpga_out_csr_writedata_7),
	.datac(!\LessThan5~1_combout ),
	.datad(!\LessThan4~4_combout ),
	.datae(!\LessThan5~0_combout ),
	.dataf(!\LessThan4~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_threshold_writedata[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_threshold_writedata[3]~3 .extended_lut = "off";
defparam \rdclk_control_slave_threshold_writedata[3]~3 .lut_mask = 64'hFF55FF75FF51FF71;
defparam \rdclk_control_slave_threshold_writedata[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_almostfull_threshold_register[3]~1 (
	.dataa(!\rdclk_control_slave_threshold_writedata[3]~3_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_almostfull_threshold_register[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_almostfull_threshold_register[3]~1 .extended_lut = "off";
defparam \rdclk_control_slave_almostfull_threshold_register[3]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdclk_control_slave_almostfull_threshold_register[3]~1 .shared_arith = "off";

dffeas \rdclk_control_slave_almostfull_threshold_register[3] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_almostfull_threshold_register[3]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always25~0_combout ),
	.q(\rdclk_control_slave_almostfull_threshold_register[3]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostfull_threshold_register[3] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostfull_threshold_register[3] .power_up = "low";

cyclonev_lcell_comb \LessThan7~2 (
	.dataa(!\rdclk_control_slave_almostfull_threshold_register[3]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~13_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan7~2 .extended_lut = "off";
defparam \LessThan7~2 .lut_mask = 64'h1111111111111111;
defparam \LessThan7~2 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_almostfull_threshold_register[2]~0 (
	.dataa(!\rdclk_control_slave_threshold_writedata[2]~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_almostfull_threshold_register[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_almostfull_threshold_register[2]~0 .extended_lut = "off";
defparam \rdclk_control_slave_almostfull_threshold_register[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdclk_control_slave_almostfull_threshold_register[2]~0 .shared_arith = "off";

dffeas \rdclk_control_slave_almostfull_threshold_register[2] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_almostfull_threshold_register[2]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always25~0_combout ),
	.q(\rdclk_control_slave_almostfull_threshold_register[2]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostfull_threshold_register[2] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostfull_threshold_register[2] .power_up = "low";

cyclonev_lcell_comb \LessThan7~3 (
	.dataa(!\rdclk_control_slave_almostfull_threshold_register[0]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~1_sumout ),
	.datac(!\rdclk_control_slave_almostfull_threshold_register[1]~q ),
	.datad(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~5_sumout ),
	.datae(!\rdclk_control_slave_almostfull_threshold_register[2]~q ),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~9_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan7~3 .extended_lut = "off";
defparam \LessThan7~3 .lut_mask = 64'h4F044F044F040000;
defparam \LessThan7~3 .shared_arith = "off";

cyclonev_lcell_comb \LessThan7~4 (
	.dataa(!\rdclk_control_slave_almostfull_threshold_register[2]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~9_sumout ),
	.datac(!\rdclk_control_slave_almostfull_threshold_register[3]~q ),
	.datad(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~13_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan7~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan7~4 .extended_lut = "off";
defparam \LessThan7~4 .lut_mask = 64'hF880F880F880F880;
defparam \LessThan7~4 .shared_arith = "off";

cyclonev_lcell_comb \LessThan7~5 (
	.dataa(!\rdclk_control_slave_almostfull_threshold_register[4]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~17_sumout ),
	.datac(!\LessThan7~1_combout ),
	.datad(!\LessThan7~2_combout ),
	.datae(!\LessThan7~3_combout ),
	.dataf(!\LessThan7~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan7~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan7~5 .extended_lut = "off";
defparam \LessThan7~5 .lut_mask = 64'h08080E080E0E0E0E;
defparam \LessThan7~5 .shared_arith = "off";

cyclonev_lcell_comb \LessThan7~6 (
	.dataa(!\rdclk_control_slave_almostfull_threshold_register[6]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~25_sumout ),
	.datac(!\rdclk_control_slave_almostfull_threshold_register[7]~q ),
	.datad(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~29_sumout ),
	.datae(!\LessThan7~0_combout ),
	.dataf(!\LessThan7~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan7~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan7~6 .extended_lut = "off";
defparam \LessThan7~6 .lut_mask = 64'hF880FEE0FEE0FEE0;
defparam \LessThan7~6 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_status_almostfull_q~0 (
	.dataa(!\LessThan7~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_status_almostfull_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_status_almostfull_q~0 .extended_lut = "off";
defparam \rdclk_control_slave_status_almostfull_q~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdclk_control_slave_status_almostfull_q~0 .shared_arith = "off";

dffeas rdclk_control_slave_status_almostfull_q(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_status_almostfull_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_status_almostfull_q~q ),
	.prn(vcc));
defparam rdclk_control_slave_status_almostfull_q.is_wysiwyg = "true";
defparam rdclk_control_slave_status_almostfull_q.power_up = "low";

cyclonev_lcell_comb \LessThan7~7 (
	.dataa(!\rdclk_control_slave_almostfull_threshold_register[2]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~9_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan7~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan7~7 .extended_lut = "off";
defparam \LessThan7~7 .lut_mask = 64'h8888888888888888;
defparam \LessThan7~7 .shared_arith = "off";

cyclonev_lcell_comb \LessThan7~8 (
	.dataa(!\rdclk_control_slave_almostfull_threshold_register[3]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~13_sumout ),
	.datac(!\rdclk_control_slave_almostfull_threshold_register[4]~q ),
	.datad(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~17_sumout ),
	.datae(!\LessThan7~3_combout ),
	.dataf(!\LessThan7~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan7~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan7~8 .extended_lut = "off";
defparam \LessThan7~8 .lut_mask = 64'h077F011F011F011F;
defparam \LessThan7~8 .shared_arith = "off";

cyclonev_lcell_comb \LessThan7~9 (
	.dataa(!\rdclk_control_slave_almostfull_threshold_register[5]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~21_sumout ),
	.datac(!\rdclk_control_slave_almostfull_threshold_register[6]~q ),
	.datad(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~25_sumout ),
	.datae(!\LessThan7~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan7~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan7~9 .extended_lut = "off";
defparam \LessThan7~9 .lut_mask = 64'hFEE0F880FEE0F880;
defparam \LessThan7~9 .shared_arith = "off";

cyclonev_lcell_comb \always30~0 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!fifo_hps_to_fpga_out_csr_write),
	.datae(!rdclk_control_slave_writedata[2]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always30~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always30~0 .extended_lut = "off";
defparam \always30~0 .lut_mask = 64'h0000000800000008;
defparam \always30~0 .shared_arith = "off";

dffeas rdclk_control_slave_almostfull_n_reg(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\LessThan7~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_almostfull_n_reg~q ),
	.prn(vcc));
defparam rdclk_control_slave_almostfull_n_reg.is_wysiwyg = "true";
defparam rdclk_control_slave_almostfull_n_reg.power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_event_almostfull_q~0 (
	.dataa(!\rdclk_control_slave_event_almostfull_q~q ),
	.datab(!\rdclk_control_slave_almostfull_threshold_register[7]~q ),
	.datac(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~29_sumout ),
	.datad(!\LessThan7~9_combout ),
	.datae(!\always30~0_combout ),
	.dataf(!\rdclk_control_slave_almostfull_n_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_event_almostfull_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_event_almostfull_q~0 .extended_lut = "off";
defparam \rdclk_control_slave_event_almostfull_q~0 .lut_mask = 64'h555500007F570000;
defparam \rdclk_control_slave_event_almostfull_q~0 .shared_arith = "off";

dffeas rdclk_control_slave_event_almostfull_q(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_event_almostfull_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_event_almostfull_q~q ),
	.prn(vcc));
defparam rdclk_control_slave_event_almostfull_q.is_wysiwyg = "true";
defparam rdclk_control_slave_event_almostfull_q.power_up = "low";

dffeas \rdclk_control_slave_ienable_register[2] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(rdclk_control_slave_writedata[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always26~0_combout ),
	.q(\rdclk_control_slave_ienable_register[2]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_ienable_register[2] .is_wysiwyg = "true";
defparam \rdclk_control_slave_ienable_register[2] .power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[2]~2 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!\rdclk_control_slave_status_almostfull_q~q ),
	.datae(!\rdclk_control_slave_event_almostfull_q~q ),
	.dataf(!\rdclk_control_slave_ienable_register[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[2]~2 .extended_lut = "off";
defparam \rdclk_control_slave_read_mux[2]~2 .lut_mask = 64'h0020082802220A2A;
defparam \rdclk_control_slave_read_mux[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[2]~20 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_1),
	.datab(!fifo_hps_to_fpga_out_csr_address_2),
	.datac(!\rdclk_control_slave_almostempty_threshold_register[2]~q ),
	.datad(!\rdclk_control_slave_read_mux[2]~2_combout ),
	.datae(!fifo_hps_to_fpga_out_csr_address_0),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~9_sumout ),
	.datag(!\rdclk_control_slave_almostfull_threshold_register[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[2]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[2]~20 .extended_lut = "on";
defparam \rdclk_control_slave_read_mux[2]~20 .lut_mask = 64'h20FF02FFB9FF13FF;
defparam \rdclk_control_slave_read_mux[2]~20 .shared_arith = "off";

dffeas \rdclk_control_slave_almostempty_threshold_register[3] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_threshold_writedata[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always24~0_combout ),
	.q(\rdclk_control_slave_almostempty_threshold_register[3]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostempty_threshold_register[3] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostempty_threshold_register[3] .power_up = "low";

dffeas \rdclk_control_slave_almostempty_threshold_register[6] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_threshold_writedata[6]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always24~0_combout ),
	.q(\rdclk_control_slave_almostempty_threshold_register[6]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostempty_threshold_register[6] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostempty_threshold_register[6] .power_up = "low";

dffeas \rdclk_control_slave_almostempty_threshold_register[7] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_threshold_writedata[7]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always24~0_combout ),
	.q(\rdclk_control_slave_almostempty_threshold_register[7]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostempty_threshold_register[7] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostempty_threshold_register[7] .power_up = "low";

dffeas \rdclk_control_slave_almostempty_threshold_register[5] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_threshold_writedata[5]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always24~0_combout ),
	.q(\rdclk_control_slave_almostempty_threshold_register[5]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostempty_threshold_register[5] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostempty_threshold_register[5] .power_up = "low";

cyclonev_lcell_comb \LessThan6~0 (
	.dataa(!\rdclk_control_slave_almostempty_threshold_register[5]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~21_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan6~0 .extended_lut = "off";
defparam \LessThan6~0 .lut_mask = 64'h2222222222222222;
defparam \LessThan6~0 .shared_arith = "off";

dffeas \rdclk_control_slave_almostempty_threshold_register[4] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_threshold_writedata[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always24~0_combout ),
	.q(\rdclk_control_slave_almostempty_threshold_register[4]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_almostempty_threshold_register[4] .is_wysiwyg = "true";
defparam \rdclk_control_slave_almostempty_threshold_register[4] .power_up = "low";

cyclonev_lcell_comb \LessThan6~1 (
	.dataa(!\rdclk_control_slave_almostempty_threshold_register[5]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~21_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan6~1 .extended_lut = "off";
defparam \LessThan6~1 .lut_mask = 64'h6666666666666666;
defparam \LessThan6~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan6~2 (
	.dataa(!\rdclk_control_slave_almostempty_threshold_register[3]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~13_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan6~2 .extended_lut = "off";
defparam \LessThan6~2 .lut_mask = 64'h4444444444444444;
defparam \LessThan6~2 .shared_arith = "off";

cyclonev_lcell_comb \LessThan6~3 (
	.dataa(!\rdclk_control_slave_almostempty_threshold_register[0]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~1_sumout ),
	.datac(!\rdclk_control_slave_almostempty_threshold_register[1]~q ),
	.datad(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~5_sumout ),
	.datae(!\rdclk_control_slave_almostempty_threshold_register[2]~q ),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~9_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan6~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan6~3 .extended_lut = "off";
defparam \LessThan6~3 .lut_mask = 64'h10F1000010F110F1;
defparam \LessThan6~3 .shared_arith = "off";

cyclonev_lcell_comb \LessThan6~4 (
	.dataa(!\rdclk_control_slave_almostempty_threshold_register[2]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~9_sumout ),
	.datac(!\rdclk_control_slave_almostempty_threshold_register[3]~q ),
	.datad(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~13_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan6~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan6~4 .extended_lut = "off";
defparam \LessThan6~4 .lut_mask = 64'h20F220F220F220F2;
defparam \LessThan6~4 .shared_arith = "off";

cyclonev_lcell_comb \LessThan6~5 (
	.dataa(!\rdclk_control_slave_almostempty_threshold_register[4]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~17_sumout ),
	.datac(!\LessThan6~1_combout ),
	.datad(!\LessThan6~2_combout ),
	.datae(!\LessThan6~3_combout ),
	.dataf(!\LessThan6~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan6~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan6~5 .extended_lut = "off";
defparam \LessThan6~5 .lut_mask = 64'h2020B020B0B0B0B0;
defparam \LessThan6~5 .shared_arith = "off";

cyclonev_lcell_comb \LessThan6~6 (
	.dataa(!\rdclk_control_slave_almostempty_threshold_register[6]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~25_sumout ),
	.datac(!\rdclk_control_slave_almostempty_threshold_register[7]~q ),
	.datad(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~29_sumout ),
	.datae(!\LessThan6~0_combout ),
	.dataf(!\LessThan6~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan6~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan6~6 .extended_lut = "off";
defparam \LessThan6~6 .lut_mask = 64'h20F2B0FBB0FBB0FB;
defparam \LessThan6~6 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_status_almostempty_q~0 (
	.dataa(!\LessThan6~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_status_almostempty_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_status_almostempty_q~0 .extended_lut = "off";
defparam \rdclk_control_slave_status_almostempty_q~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdclk_control_slave_status_almostempty_q~0 .shared_arith = "off";

dffeas rdclk_control_slave_status_almostempty_q(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_status_almostempty_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_status_almostempty_q~q ),
	.prn(vcc));
defparam rdclk_control_slave_status_almostempty_q.is_wysiwyg = "true";
defparam rdclk_control_slave_status_almostempty_q.power_up = "low";

cyclonev_lcell_comb \LessThan6~7 (
	.dataa(!\rdclk_control_slave_almostempty_threshold_register[2]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~9_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan6~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan6~7 .extended_lut = "off";
defparam \LessThan6~7 .lut_mask = 64'h2222222222222222;
defparam \LessThan6~7 .shared_arith = "off";

cyclonev_lcell_comb \LessThan6~8 (
	.dataa(!\rdclk_control_slave_almostempty_threshold_register[3]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~13_sumout ),
	.datac(!\rdclk_control_slave_almostempty_threshold_register[4]~q ),
	.datad(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~17_sumout ),
	.datae(!\LessThan6~3_combout ),
	.dataf(!\LessThan6~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan6~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan6~8 .extended_lut = "off";
defparam \LessThan6~8 .lut_mask = 64'hDF0D4F044F044F04;
defparam \LessThan6~8 .shared_arith = "off";

cyclonev_lcell_comb \LessThan6~9 (
	.dataa(!\rdclk_control_slave_almostempty_threshold_register[5]~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~21_sumout ),
	.datac(!\rdclk_control_slave_almostempty_threshold_register[6]~q ),
	.datad(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~25_sumout ),
	.datae(!\LessThan6~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan6~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan6~9 .extended_lut = "off";
defparam \LessThan6~9 .lut_mask = 64'hB0FB20F2B0FB20F2;
defparam \LessThan6~9 .shared_arith = "off";

cyclonev_lcell_comb \always29~0 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!fifo_hps_to_fpga_out_csr_write),
	.datae(!rdclk_control_slave_writedata[3]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always29~0 .extended_lut = "off";
defparam \always29~0 .lut_mask = 64'h0000000800000008;
defparam \always29~0 .shared_arith = "off";

dffeas rdclk_control_slave_almostempty_n_reg(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\LessThan6~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_almostempty_n_reg~q ),
	.prn(vcc));
defparam rdclk_control_slave_almostempty_n_reg.is_wysiwyg = "true";
defparam rdclk_control_slave_almostempty_n_reg.power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_event_almostempty_q~0 (
	.dataa(!\rdclk_control_slave_event_almostempty_q~q ),
	.datab(!\rdclk_control_slave_almostempty_threshold_register[7]~q ),
	.datac(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~29_sumout ),
	.datad(!\LessThan6~9_combout ),
	.datae(!\always29~0_combout ),
	.dataf(!\rdclk_control_slave_almostempty_n_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_event_almostempty_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_event_almostempty_q~0 .extended_lut = "off";
defparam \rdclk_control_slave_event_almostempty_q~0 .lut_mask = 64'h55550000F7750000;
defparam \rdclk_control_slave_event_almostempty_q~0 .shared_arith = "off";

dffeas rdclk_control_slave_event_almostempty_q(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_event_almostempty_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_event_almostempty_q~q ),
	.prn(vcc));
defparam rdclk_control_slave_event_almostempty_q.is_wysiwyg = "true";
defparam rdclk_control_slave_event_almostempty_q.power_up = "low";

dffeas \rdclk_control_slave_ienable_register[3] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(rdclk_control_slave_writedata[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always26~0_combout ),
	.q(\rdclk_control_slave_ienable_register[3]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_ienable_register[3] .is_wysiwyg = "true";
defparam \rdclk_control_slave_ienable_register[3] .power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[3]~3 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!\rdclk_control_slave_status_almostempty_q~q ),
	.datae(!\rdclk_control_slave_event_almostempty_q~q ),
	.dataf(!\rdclk_control_slave_ienable_register[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[3]~3 .extended_lut = "off";
defparam \rdclk_control_slave_read_mux[3]~3 .lut_mask = 64'h0020082802220A2A;
defparam \rdclk_control_slave_read_mux[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[3]~16 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_1),
	.datab(!fifo_hps_to_fpga_out_csr_address_2),
	.datac(!\rdclk_control_slave_almostempty_threshold_register[3]~q ),
	.datad(!\rdclk_control_slave_read_mux[3]~3_combout ),
	.datae(!fifo_hps_to_fpga_out_csr_address_0),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~13_sumout ),
	.datag(!\rdclk_control_slave_almostfull_threshold_register[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[3]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[3]~16 .extended_lut = "on";
defparam \rdclk_control_slave_read_mux[3]~16 .lut_mask = 64'h20FF02FFB9FF13FF;
defparam \rdclk_control_slave_read_mux[3]~16 .shared_arith = "off";

cyclonev_lcell_comb rdclk_control_slave_status_overflow_signal(
	.dataa(!\the_dcfifo|dual_clock_fifo|auto_generated|rdfull_eq_comp|aneb_result_wire[0]~3_combout ),
	.datab(!\the_dcfifo|rdfull~0_combout ),
	.datac(!\the_dcfifo|rdfull~1_combout ),
	.datad(!\wrdreq_sync_i|dreg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_status_overflow_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam rdclk_control_slave_status_overflow_signal.extended_lut = "off";
defparam rdclk_control_slave_status_overflow_signal.lut_mask = 64'h0057005700570057;
defparam rdclk_control_slave_status_overflow_signal.shared_arith = "off";

dffeas rdclk_control_slave_status_overflow_q(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_status_overflow_signal~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_status_overflow_q~q ),
	.prn(vcc));
defparam rdclk_control_slave_status_overflow_q.is_wysiwyg = "true";
defparam rdclk_control_slave_status_overflow_q.power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_event_overflow_q~0 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!fifo_hps_to_fpga_out_csr_write),
	.datae(!rdclk_control_slave_writedata[4]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_event_overflow_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_event_overflow_q~0 .extended_lut = "off";
defparam \rdclk_control_slave_event_overflow_q~0 .lut_mask = 64'h0000000800000008;
defparam \rdclk_control_slave_event_overflow_q~0 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_event_overflow_q~1 (
	.dataa(!\rdclk_control_slave_event_overflow_q~q ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|rdfull_eq_comp|aneb_result_wire[0]~3_combout ),
	.datac(!\the_dcfifo|rdfull~0_combout ),
	.datad(!\the_dcfifo|rdfull~1_combout ),
	.datae(!\wrdreq_sync_i|dreg[2]~q ),
	.dataf(!\rdclk_control_slave_event_overflow_q~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_event_overflow_q~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_event_overflow_q~1 .extended_lut = "off";
defparam \rdclk_control_slave_event_overflow_q~1 .lut_mask = 64'h5555777F00000000;
defparam \rdclk_control_slave_event_overflow_q~1 .shared_arith = "off";

dffeas rdclk_control_slave_event_overflow_q(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_event_overflow_q~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_event_overflow_q~q ),
	.prn(vcc));
defparam rdclk_control_slave_event_overflow_q.is_wysiwyg = "true";
defparam rdclk_control_slave_event_overflow_q.power_up = "low";

dffeas \rdclk_control_slave_ienable_register[4] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(rdclk_control_slave_writedata[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always26~0_combout ),
	.q(\rdclk_control_slave_ienable_register[4]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_ienable_register[4] .is_wysiwyg = "true";
defparam \rdclk_control_slave_ienable_register[4] .power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[4]~4 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!\rdclk_control_slave_status_overflow_q~q ),
	.datae(!\rdclk_control_slave_event_overflow_q~q ),
	.dataf(!\rdclk_control_slave_ienable_register[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[4]~4 .extended_lut = "off";
defparam \rdclk_control_slave_read_mux[4]~4 .lut_mask = 64'h0020082802220A2A;
defparam \rdclk_control_slave_read_mux[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[4]~12 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_1),
	.datab(!fifo_hps_to_fpga_out_csr_address_2),
	.datac(!\rdclk_control_slave_almostempty_threshold_register[4]~q ),
	.datad(!\rdclk_control_slave_read_mux[4]~4_combout ),
	.datae(!fifo_hps_to_fpga_out_csr_address_0),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~17_sumout ),
	.datag(!\rdclk_control_slave_almostfull_threshold_register[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[4]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[4]~12 .extended_lut = "on";
defparam \rdclk_control_slave_read_mux[4]~12 .lut_mask = 64'h20FF02FFB9FF13FF;
defparam \rdclk_control_slave_read_mux[4]~12 .shared_arith = "off";

cyclonev_lcell_comb rdclk_control_slave_status_underflow_signal(
	.dataa(!\the_dcfifo|dual_clock_fifo|auto_generated|rdempty_eq_comp|data_wire[2]~0_combout ),
	.datab(!fifo_hps_to_fpga_out_read),
	.datac(!\the_dcfifo|dual_clock_fifo|auto_generated|rdfull_eq_comp|aneb_result_wire[0]~0_combout ),
	.datad(!\the_dcfifo|dual_clock_fifo|auto_generated|rdfull_eq_comp|aneb_result_wire[0]~1_combout ),
	.datae(!\the_dcfifo|dual_clock_fifo|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_status_underflow_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam rdclk_control_slave_status_underflow_signal.extended_lut = "off";
defparam rdclk_control_slave_status_underflow_signal.lut_mask = 64'h0000000200000002;
defparam rdclk_control_slave_status_underflow_signal.shared_arith = "off";

dffeas rdclk_control_slave_status_underflow_q(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_status_underflow_signal~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_status_underflow_q~q ),
	.prn(vcc));
defparam rdclk_control_slave_status_underflow_q.is_wysiwyg = "true";
defparam rdclk_control_slave_status_underflow_q.power_up = "low";

cyclonev_lcell_comb \always29~1 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!fifo_hps_to_fpga_out_csr_write),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always29~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always29~1 .extended_lut = "off";
defparam \always29~1 .lut_mask = 64'h0008000800080008;
defparam \always29~1 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_event_underflow_q~0 (
	.dataa(!\rdclk_control_slave_event_underflow_q~q ),
	.datab(!\always29~1_combout ),
	.datac(!rdclk_control_slave_writedata[5]),
	.datad(!\rdclk_control_slave_status_underflow_signal~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_event_underflow_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_event_underflow_q~0 .extended_lut = "off";
defparam \rdclk_control_slave_event_underflow_q~0 .lut_mask = 64'h54FC54FC54FC54FC;
defparam \rdclk_control_slave_event_underflow_q~0 .shared_arith = "off";

dffeas rdclk_control_slave_event_underflow_q(
	.clk(clock_bridge_0_in_clk_clk),
	.d(\rdclk_control_slave_event_underflow_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdclk_control_slave_event_underflow_q~q ),
	.prn(vcc));
defparam rdclk_control_slave_event_underflow_q.is_wysiwyg = "true";
defparam rdclk_control_slave_event_underflow_q.power_up = "low";

dffeas \rdclk_control_slave_ienable_register[5] (
	.clk(clock_bridge_0_in_clk_clk),
	.d(rdclk_control_slave_writedata[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always26~0_combout ),
	.q(\rdclk_control_slave_ienable_register[5]~q ),
	.prn(vcc));
defparam \rdclk_control_slave_ienable_register[5] .is_wysiwyg = "true";
defparam \rdclk_control_slave_ienable_register[5] .power_up = "low";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[5]~5 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!\rdclk_control_slave_status_underflow_q~q ),
	.datae(!\rdclk_control_slave_event_underflow_q~q ),
	.dataf(!\rdclk_control_slave_ienable_register[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[5]~5 .extended_lut = "off";
defparam \rdclk_control_slave_read_mux[5]~5 .lut_mask = 64'h0020082802220A2A;
defparam \rdclk_control_slave_read_mux[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[5]~8 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_1),
	.datab(!fifo_hps_to_fpga_out_csr_address_2),
	.datac(!\rdclk_control_slave_almostempty_threshold_register[5]~q ),
	.datad(!\rdclk_control_slave_read_mux[5]~5_combout ),
	.datae(!fifo_hps_to_fpga_out_csr_address_0),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~21_sumout ),
	.datag(!\rdclk_control_slave_almostfull_threshold_register[5]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[5]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[5]~8 .extended_lut = "on";
defparam \rdclk_control_slave_read_mux[5]~8 .lut_mask = 64'h20FF02FFB9FF13FF;
defparam \rdclk_control_slave_read_mux[5]~8 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[6]~6 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!\rdclk_control_slave_almostfull_threshold_register[6]~q ),
	.datae(!\rdclk_control_slave_almostempty_threshold_register[6]~q ),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~25_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[6]~6 .extended_lut = "off";
defparam \rdclk_control_slave_read_mux[6]~6 .lut_mask = 64'h40005010C585D595;
defparam \rdclk_control_slave_read_mux[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \rdclk_control_slave_read_mux[7]~7 (
	.dataa(!fifo_hps_to_fpga_out_csr_address_2),
	.datab(!fifo_hps_to_fpga_out_csr_address_0),
	.datac(!fifo_hps_to_fpga_out_csr_address_1),
	.datad(!\rdclk_control_slave_almostfull_threshold_register[7]~q ),
	.datae(!\rdclk_control_slave_almostempty_threshold_register[7]~q ),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_1~29_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdclk_control_slave_read_mux[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdclk_control_slave_read_mux[7]~7 .extended_lut = "off";
defparam \rdclk_control_slave_read_mux[7]~7 .lut_mask = 64'h40005010C585D595;
defparam \rdclk_control_slave_read_mux[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!in_data_reg_131),
	.datab(!in_data_reg_121),
	.datac(!in_data_reg_111),
	.datad(!in_data_reg_101),
	.datae(!in_data_reg_91),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8000000080000000;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!in_data_reg_191),
	.datab(!in_data_reg_181),
	.datac(!in_data_reg_171),
	.datad(!in_data_reg_161),
	.datae(!in_data_reg_151),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h8000000080000000;
defparam \LessThan0~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~2 (
	.dataa(!in_data_reg_311),
	.datab(!in_data_reg_301),
	.datac(!in_data_reg_291),
	.datad(!in_data_reg_281),
	.datae(!in_data_reg_271),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~2 .extended_lut = "off";
defparam \LessThan0~2 .lut_mask = 64'h8000000080000000;
defparam \LessThan0~2 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~3 (
	.dataa(!in_data_reg_251),
	.datab(!in_data_reg_241),
	.datac(!in_data_reg_231),
	.datad(!in_data_reg_221),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~3 .extended_lut = "off";
defparam \LessThan0~3 .lut_mask = 64'h8000800080008000;
defparam \LessThan0~3 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~4 (
	.dataa(!in_data_reg_261),
	.datab(!in_data_reg_211),
	.datac(!in_data_reg_201),
	.datad(!\LessThan0~2_combout ),
	.datae(!\LessThan0~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~4 .extended_lut = "off";
defparam \LessThan0~4 .lut_mask = 64'h0000008000000080;
defparam \LessThan0~4 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~5 (
	.dataa(!in_data_reg_141),
	.datab(!in_data_reg_81),
	.datac(!\LessThan0~0_combout ),
	.datad(!\LessThan0~1_combout ),
	.datae(!\LessThan0~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~5 .extended_lut = "off";
defparam \LessThan0~5 .lut_mask = 64'h0000000800000008;
defparam \LessThan0~5 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~0 (
	.dataa(!in_data_reg_71),
	.datab(!in_data_reg_61),
	.datac(!wrclk_control_slave_writedata[5]),
	.datad(!wrclk_control_slave_writedata[4]),
	.datae(!wrclk_control_slave_writedata[3]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~0 .extended_lut = "off";
defparam \LessThan1~0 .lut_mask = 64'h0000000100000001;
defparam \LessThan1~0 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_threshold_writedata~0 (
	.dataa(!wrclk_control_slave_writedata[0]),
	.datab(!wrclk_control_slave_writedata[2]),
	.datac(!wrclk_control_slave_writedata[1]),
	.datad(!\LessThan0~5_combout ),
	.datae(!\LessThan1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_threshold_writedata~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_threshold_writedata~0 .extended_lut = "off";
defparam \wrclk_control_slave_threshold_writedata~0 .lut_mask = 64'h00FF00EC00FF00EC;
defparam \wrclk_control_slave_threshold_writedata~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~6 (
	.dataa(!in_data_reg_71),
	.datab(!in_data_reg_61),
	.datac(!wrclk_control_slave_writedata[5]),
	.datad(!wrclk_control_slave_writedata[4]),
	.datae(!wrclk_control_slave_writedata[3]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~6 .extended_lut = "off";
defparam \LessThan0~6 .lut_mask = 64'h8000000080000000;
defparam \LessThan0~6 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~7 (
	.dataa(!wrclk_control_slave_writedata[0]),
	.datab(!wrclk_control_slave_writedata[2]),
	.datac(!wrclk_control_slave_writedata[1]),
	.datad(!\LessThan0~5_combout ),
	.datae(!\LessThan0~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~7 .extended_lut = "off";
defparam \LessThan0~7 .lut_mask = 64'h0000008000000080;
defparam \LessThan0~7 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_threshold_writedata[0]~1 (
	.dataa(!wrclk_control_slave_writedata[0]),
	.datab(!\wrclk_control_slave_threshold_writedata~0_combout ),
	.datac(!\LessThan0~7_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_threshold_writedata[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_threshold_writedata[0]~1 .extended_lut = "off";
defparam \wrclk_control_slave_threshold_writedata[0]~1 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \wrclk_control_slave_threshold_writedata[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_almostempty_threshold_register[0]~0 (
	.dataa(!\wrclk_control_slave_threshold_writedata[0]~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_almostempty_threshold_register[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_almostempty_threshold_register[0]~0 .extended_lut = "off";
defparam \wrclk_control_slave_almostempty_threshold_register[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wrclk_control_slave_almostempty_threshold_register[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \always4~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!m0_write1),
	.datac(!wait_latency_counter_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'h2020202020202020;
defparam \always4~0 .shared_arith = "off";

cyclonev_lcell_comb \always4~1 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!\always4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~1 .extended_lut = "off";
defparam \always4~1 .lut_mask = 64'h0010001000100010;
defparam \always4~1 .shared_arith = "off";

dffeas \wrclk_control_slave_almostempty_threshold_register[0] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_almostempty_threshold_register[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\wrclk_control_slave_almostempty_threshold_register[0]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostempty_threshold_register[0] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostempty_threshold_register[0] .power_up = "low";

dffeas wrclk_control_slave_status_full_q(
	.clk(outclk_wire_0),
	.d(\the_dcfifo|wrfull~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_status_full_q~q ),
	.prn(vcc));
defparam wrclk_control_slave_status_full_q.is_wysiwyg = "true";
defparam wrclk_control_slave_status_full_q.power_up = "low";

cyclonev_lcell_comb \always7~0 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!\always4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always7~0 .extended_lut = "off";
defparam \always7~0 .lut_mask = 64'h0008000800080008;
defparam \always7~0 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_full_n_reg~0 (
	.dataa(!\the_dcfifo|wrfull~7_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_full_n_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_full_n_reg~0 .extended_lut = "off";
defparam \wrclk_control_slave_full_n_reg~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wrclk_control_slave_full_n_reg~0 .shared_arith = "off";

dffeas wrclk_control_slave_full_n_reg(
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_full_n_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_full_n_reg~q ),
	.prn(vcc));
defparam wrclk_control_slave_full_n_reg.is_wysiwyg = "true";
defparam wrclk_control_slave_full_n_reg.power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_event_full_q~0 (
	.dataa(!\the_dcfifo|wrfull~7_combout ),
	.datab(!\wrclk_control_slave_event_full_q~q ),
	.datac(!wrclk_control_slave_writedata[0]),
	.datad(!\always7~0_combout ),
	.datae(!\wrclk_control_slave_full_n_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_event_full_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_event_full_q~0 .extended_lut = "off";
defparam \wrclk_control_slave_event_full_q~0 .lut_mask = 64'h3330777033307770;
defparam \wrclk_control_slave_event_full_q~0 .shared_arith = "off";

dffeas wrclk_control_slave_event_full_q(
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_event_full_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_event_full_q~q ),
	.prn(vcc));
defparam wrclk_control_slave_event_full_q.is_wysiwyg = "true";
defparam wrclk_control_slave_event_full_q.power_up = "low";

cyclonev_lcell_comb \always6~0 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!\always4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~0 .extended_lut = "off";
defparam \always6~0 .lut_mask = 64'h0004000400040004;
defparam \always6~0 .shared_arith = "off";

dffeas \wrclk_control_slave_ienable_register[0] (
	.clk(outclk_wire_0),
	.d(wrclk_control_slave_writedata[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\wrclk_control_slave_ienable_register[0]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_ienable_register[0] .is_wysiwyg = "true";
defparam \wrclk_control_slave_ienable_register[0] .power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[0]~0 (
	.dataa(!\wrclk_control_slave_status_full_q~q ),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\wrclk_control_slave_event_full_q~q ),
	.dataf(!\wrclk_control_slave_ienable_register[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[0]~0 .extended_lut = "off";
defparam \wrclk_control_slave_read_mux[0]~0 .lut_mask = 64'h100010C0103010F0;
defparam \wrclk_control_slave_read_mux[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \always5~0 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!\always4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always5~0 .extended_lut = "off";
defparam \always5~0 .lut_mask = 64'h0020002000200020;
defparam \always5~0 .shared_arith = "off";

dffeas \wrclk_control_slave_almostfull_threshold_register[0] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_threshold_writedata[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\wrclk_control_slave_almostfull_threshold_register[0]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostfull_threshold_register[0] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostfull_threshold_register[0] .power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[0]~28 (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!\wrclk_control_slave_almostempty_threshold_register[0]~q ),
	.datad(!\wrclk_control_slave_read_mux[0]~0_combout ),
	.datae(!int_nxt_addr_reg_dly_2),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~17_sumout ),
	.datag(!\wrclk_control_slave_almostfull_threshold_register[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[0]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[0]~28 .extended_lut = "on";
defparam \wrclk_control_slave_read_mux[0]~28 .lut_mask = 64'h02FF20FF9BFF31FF;
defparam \wrclk_control_slave_read_mux[0]~28 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_threshold_writedata[1]~2 (
	.dataa(!wrclk_control_slave_writedata[1]),
	.datab(!\wrclk_control_slave_threshold_writedata~0_combout ),
	.datac(!\LessThan0~7_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_threshold_writedata[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_threshold_writedata[1]~2 .extended_lut = "off";
defparam \wrclk_control_slave_threshold_writedata[1]~2 .lut_mask = 64'h1010101010101010;
defparam \wrclk_control_slave_threshold_writedata[1]~2 .shared_arith = "off";

dffeas \wrclk_control_slave_almostempty_threshold_register[1] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_threshold_writedata[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\wrclk_control_slave_almostempty_threshold_register[1]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostempty_threshold_register[1] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostempty_threshold_register[1] .power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_status_empty_q~0 (
	.dataa(!\the_dcfifo|dual_clock_fifo|auto_generated|wrempty_eq_comp|aneb_result_wire[0]~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_status_empty_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_status_empty_q~0 .extended_lut = "off";
defparam \wrclk_control_slave_status_empty_q~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wrclk_control_slave_status_empty_q~0 .shared_arith = "off";

dffeas wrclk_control_slave_status_empty_q(
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_status_empty_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_status_empty_q~q ),
	.prn(vcc));
defparam wrclk_control_slave_status_empty_q.is_wysiwyg = "true";
defparam wrclk_control_slave_status_empty_q.power_up = "low";

dffeas wrclk_control_slave_empty_n_reg(
	.clk(outclk_wire_0),
	.d(\the_dcfifo|dual_clock_fifo|auto_generated|wrempty_eq_comp|aneb_result_wire[0]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_empty_n_reg~q ),
	.prn(vcc));
defparam wrclk_control_slave_empty_n_reg.is_wysiwyg = "true";
defparam wrclk_control_slave_empty_n_reg.power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_event_empty_q~0 (
	.dataa(!\wrclk_control_slave_event_empty_q~q ),
	.datab(!\always7~0_combout ),
	.datac(!wrclk_control_slave_writedata[1]),
	.datad(!\wrclk_control_slave_empty_n_reg~q ),
	.datae(!\the_dcfifo|dual_clock_fifo|auto_generated|wrempty_eq_comp|aneb_result_wire[0]~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_event_empty_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_event_empty_q~0 .extended_lut = "off";
defparam \wrclk_control_slave_event_empty_q~0 .lut_mask = 64'h54FC545454FC5454;
defparam \wrclk_control_slave_event_empty_q~0 .shared_arith = "off";

dffeas wrclk_control_slave_event_empty_q(
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_event_empty_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_event_empty_q~q ),
	.prn(vcc));
defparam wrclk_control_slave_event_empty_q.is_wysiwyg = "true";
defparam wrclk_control_slave_event_empty_q.power_up = "low";

dffeas \wrclk_control_slave_ienable_register[1] (
	.clk(outclk_wire_0),
	.d(wrclk_control_slave_writedata[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\wrclk_control_slave_ienable_register[1]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_ienable_register[1] .is_wysiwyg = "true";
defparam \wrclk_control_slave_ienable_register[1] .power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[1]~1 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!\wrclk_control_slave_status_empty_q~q ),
	.datae(!\wrclk_control_slave_event_empty_q~q ),
	.dataf(!\wrclk_control_slave_ienable_register[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[1]~1 .extended_lut = "off";
defparam \wrclk_control_slave_read_mux[1]~1 .lut_mask = 64'h0040084804440C4C;
defparam \wrclk_control_slave_read_mux[1]~1 .shared_arith = "off";

dffeas \wrclk_control_slave_almostfull_threshold_register[1] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_threshold_writedata[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\wrclk_control_slave_almostfull_threshold_register[1]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostfull_threshold_register[1] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostfull_threshold_register[1] .power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[1]~24 (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!\wrclk_control_slave_almostempty_threshold_register[1]~q ),
	.datad(!\wrclk_control_slave_read_mux[1]~1_combout ),
	.datae(!int_nxt_addr_reg_dly_2),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~21_sumout ),
	.datag(!\wrclk_control_slave_almostfull_threshold_register[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[1]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[1]~24 .extended_lut = "on";
defparam \wrclk_control_slave_read_mux[1]~24 .lut_mask = 64'h02FF02FF9BFF13FF;
defparam \wrclk_control_slave_read_mux[1]~24 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_threshold_writedata[2]~3 (
	.dataa(!wrclk_control_slave_writedata[2]),
	.datab(!\wrclk_control_slave_threshold_writedata~0_combout ),
	.datac(!\LessThan0~7_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_threshold_writedata[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_threshold_writedata[2]~3 .extended_lut = "off";
defparam \wrclk_control_slave_threshold_writedata[2]~3 .lut_mask = 64'hD0D0D0D0D0D0D0D0;
defparam \wrclk_control_slave_threshold_writedata[2]~3 .shared_arith = "off";

dffeas \wrclk_control_slave_almostempty_threshold_register[2] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_threshold_writedata[2]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\wrclk_control_slave_almostempty_threshold_register[2]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostempty_threshold_register[2] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostempty_threshold_register[2] .power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_almostfull_threshold_register[2]~0 (
	.dataa(!\wrclk_control_slave_threshold_writedata[2]~3_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_almostfull_threshold_register[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_almostfull_threshold_register[2]~0 .extended_lut = "off";
defparam \wrclk_control_slave_almostfull_threshold_register[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wrclk_control_slave_almostfull_threshold_register[2]~0 .shared_arith = "off";

dffeas \wrclk_control_slave_almostfull_threshold_register[2] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_almostfull_threshold_register[2]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\wrclk_control_slave_almostfull_threshold_register[2]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostfull_threshold_register[2] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostfull_threshold_register[2] .power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_threshold_writedata[3]~4 (
	.dataa(!wrclk_control_slave_writedata[3]),
	.datab(!\wrclk_control_slave_threshold_writedata~0_combout ),
	.datac(!\LessThan0~7_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_threshold_writedata[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_threshold_writedata[3]~4 .extended_lut = "off";
defparam \wrclk_control_slave_threshold_writedata[3]~4 .lut_mask = 64'hD0D0D0D0D0D0D0D0;
defparam \wrclk_control_slave_threshold_writedata[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_almostfull_threshold_register[3]~1 (
	.dataa(!\wrclk_control_slave_threshold_writedata[3]~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_almostfull_threshold_register[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_almostfull_threshold_register[3]~1 .extended_lut = "off";
defparam \wrclk_control_slave_almostfull_threshold_register[3]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wrclk_control_slave_almostfull_threshold_register[3]~1 .shared_arith = "off";

dffeas \wrclk_control_slave_almostfull_threshold_register[3] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_almostfull_threshold_register[3]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\wrclk_control_slave_almostfull_threshold_register[3]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostfull_threshold_register[3] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostfull_threshold_register[3] .power_up = "low";

cyclonev_lcell_comb \LessThan3~0 (
	.dataa(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~17_sumout ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~21_sumout ),
	.datac(!\wrclk_control_slave_almostfull_threshold_register[0]~q ),
	.datad(!\wrclk_control_slave_almostfull_threshold_register[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~0 .extended_lut = "off";
defparam \LessThan3~0 .lut_mask = 64'h08CE08CE08CE08CE;
defparam \LessThan3~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~2 (
	.dataa(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~1_sumout ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~5_sumout ),
	.datac(!\wrclk_control_slave_almostfull_threshold_register[2]~q ),
	.datad(!\wrclk_control_slave_almostfull_threshold_register[3]~q ),
	.datae(!\LessThan3~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~2 .extended_lut = "off";
defparam \LessThan3~2 .lut_mask = 64'hEC80FEC8EC80FEC8;
defparam \LessThan3~2 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_threshold_writedata[6]~7 (
	.dataa(!in_data_reg_61),
	.datab(!\wrclk_control_slave_threshold_writedata~0_combout ),
	.datac(!\LessThan0~7_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_threshold_writedata[6]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_threshold_writedata[6]~7 .extended_lut = "off";
defparam \wrclk_control_slave_threshold_writedata[6]~7 .lut_mask = 64'hD0D0D0D0D0D0D0D0;
defparam \wrclk_control_slave_threshold_writedata[6]~7 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_almostfull_threshold_register[6]~4 (
	.dataa(!\wrclk_control_slave_threshold_writedata[6]~7_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_almostfull_threshold_register[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_almostfull_threshold_register[6]~4 .extended_lut = "off";
defparam \wrclk_control_slave_almostfull_threshold_register[6]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wrclk_control_slave_almostfull_threshold_register[6]~4 .shared_arith = "off";

dffeas \wrclk_control_slave_almostfull_threshold_register[6] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_almostfull_threshold_register[6]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\wrclk_control_slave_almostfull_threshold_register[6]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostfull_threshold_register[6] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostfull_threshold_register[6] .power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_threshold_writedata[4]~5 (
	.dataa(!wrclk_control_slave_writedata[4]),
	.datab(!\wrclk_control_slave_threshold_writedata~0_combout ),
	.datac(!\LessThan0~7_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_threshold_writedata[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_threshold_writedata[4]~5 .extended_lut = "off";
defparam \wrclk_control_slave_threshold_writedata[4]~5 .lut_mask = 64'hD0D0D0D0D0D0D0D0;
defparam \wrclk_control_slave_threshold_writedata[4]~5 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_almostfull_threshold_register[4]~2 (
	.dataa(!\wrclk_control_slave_threshold_writedata[4]~5_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_almostfull_threshold_register[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_almostfull_threshold_register[4]~2 .extended_lut = "off";
defparam \wrclk_control_slave_almostfull_threshold_register[4]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wrclk_control_slave_almostfull_threshold_register[4]~2 .shared_arith = "off";

dffeas \wrclk_control_slave_almostfull_threshold_register[4] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_almostfull_threshold_register[4]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\wrclk_control_slave_almostfull_threshold_register[4]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostfull_threshold_register[4] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostfull_threshold_register[4] .power_up = "low";

cyclonev_lcell_comb \LessThan3~3 (
	.dataa(!op_21),
	.datab(!\wrclk_control_slave_almostfull_threshold_register[6]~q ),
	.datac(!\wrclk_control_slave_almostfull_threshold_register[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~3 .extended_lut = "off";
defparam \LessThan3~3 .lut_mask = 64'hE8E8E8E8E8E8E8E8;
defparam \LessThan3~3 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_threshold_writedata[7]~8 (
	.dataa(!in_data_reg_71),
	.datab(!\wrclk_control_slave_threshold_writedata~0_combout ),
	.datac(!\LessThan0~7_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_threshold_writedata[7]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_threshold_writedata[7]~8 .extended_lut = "off";
defparam \wrclk_control_slave_threshold_writedata[7]~8 .lut_mask = 64'hD0D0D0D0D0D0D0D0;
defparam \wrclk_control_slave_threshold_writedata[7]~8 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_almostfull_threshold_register[7]~5 (
	.dataa(!\wrclk_control_slave_threshold_writedata[7]~8_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_almostfull_threshold_register[7]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_almostfull_threshold_register[7]~5 .extended_lut = "off";
defparam \wrclk_control_slave_almostfull_threshold_register[7]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wrclk_control_slave_almostfull_threshold_register[7]~5 .shared_arith = "off";

dffeas \wrclk_control_slave_almostfull_threshold_register[7] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_almostfull_threshold_register[7]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\wrclk_control_slave_almostfull_threshold_register[7]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostfull_threshold_register[7] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostfull_threshold_register[7] .power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_threshold_writedata[5]~6 (
	.dataa(!wrclk_control_slave_writedata[5]),
	.datab(!\wrclk_control_slave_threshold_writedata~0_combout ),
	.datac(!\LessThan0~7_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_threshold_writedata[5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_threshold_writedata[5]~6 .extended_lut = "off";
defparam \wrclk_control_slave_threshold_writedata[5]~6 .lut_mask = 64'hD0D0D0D0D0D0D0D0;
defparam \wrclk_control_slave_threshold_writedata[5]~6 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_almostfull_threshold_register[5]~3 (
	.dataa(!\wrclk_control_slave_threshold_writedata[5]~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_almostfull_threshold_register[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_almostfull_threshold_register[5]~3 .extended_lut = "off";
defparam \wrclk_control_slave_almostfull_threshold_register[5]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wrclk_control_slave_almostfull_threshold_register[5]~3 .shared_arith = "off";

dffeas \wrclk_control_slave_almostfull_threshold_register[5] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_almostfull_threshold_register[5]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\wrclk_control_slave_almostfull_threshold_register[5]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostfull_threshold_register[5] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostfull_threshold_register[5] .power_up = "low";

cyclonev_lcell_comb \LessThan3~4 (
	.dataa(!op_21),
	.datab(!op_22),
	.datac(!\wrclk_control_slave_almostfull_threshold_register[6]~q ),
	.datad(!\wrclk_control_slave_almostfull_threshold_register[7]~q ),
	.datae(!op_2),
	.dataf(!\wrclk_control_slave_almostfull_threshold_register[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~4 .extended_lut = "off";
defparam \LessThan3~4 .lut_mask = 64'h013701370137137F;
defparam \LessThan3~4 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~5 (
	.dataa(!op_21),
	.datab(!op_22),
	.datac(!\wrclk_control_slave_almostfull_threshold_register[6]~q ),
	.datad(!\wrclk_control_slave_almostfull_threshold_register[7]~q ),
	.datae(!op_2),
	.dataf(!\wrclk_control_slave_almostfull_threshold_register[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~5 .extended_lut = "off";
defparam \LessThan3~5 .lut_mask = 64'h0000135F135F135F;
defparam \LessThan3~5 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~1 (
	.dataa(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~9_sumout ),
	.datab(!\LessThan3~2_combout ),
	.datac(!\LessThan3~3_combout ),
	.datad(!\LessThan3~4_combout ),
	.datae(!\LessThan3~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~1 .extended_lut = "off";
defparam \LessThan3~1 .lut_mask = 64'hFF002B00FF002B00;
defparam \LessThan3~1 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_status_almostfull_q~0 (
	.dataa(!\LessThan3~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_status_almostfull_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_status_almostfull_q~0 .extended_lut = "off";
defparam \wrclk_control_slave_status_almostfull_q~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wrclk_control_slave_status_almostfull_q~0 .shared_arith = "off";

dffeas wrclk_control_slave_status_almostfull_q(
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_status_almostfull_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_status_almostfull_q~q ),
	.prn(vcc));
defparam wrclk_control_slave_status_almostfull_q.is_wysiwyg = "true";
defparam wrclk_control_slave_status_almostfull_q.power_up = "low";

dffeas wrclk_control_slave_almostfull_n_reg(
	.clk(outclk_wire_0),
	.d(\LessThan3~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_almostfull_n_reg~q ),
	.prn(vcc));
defparam wrclk_control_slave_almostfull_n_reg.is_wysiwyg = "true";
defparam wrclk_control_slave_almostfull_n_reg.power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_event_almostfull_q~0 (
	.dataa(!\wrclk_control_slave_event_almostfull_q~q ),
	.datab(!\always7~0_combout ),
	.datac(!wrclk_control_slave_writedata[2]),
	.datad(!\LessThan3~1_combout ),
	.datae(!\wrclk_control_slave_almostfull_n_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_event_almostfull_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_event_almostfull_q~0 .extended_lut = "off";
defparam \wrclk_control_slave_event_almostfull_q~0 .lut_mask = 64'h5454FC545454FC54;
defparam \wrclk_control_slave_event_almostfull_q~0 .shared_arith = "off";

dffeas wrclk_control_slave_event_almostfull_q(
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_event_almostfull_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_event_almostfull_q~q ),
	.prn(vcc));
defparam wrclk_control_slave_event_almostfull_q.is_wysiwyg = "true";
defparam wrclk_control_slave_event_almostfull_q.power_up = "low";

dffeas \wrclk_control_slave_ienable_register[2] (
	.clk(outclk_wire_0),
	.d(wrclk_control_slave_writedata[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\wrclk_control_slave_ienable_register[2]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_ienable_register[2] .is_wysiwyg = "true";
defparam \wrclk_control_slave_ienable_register[2] .power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[2]~2 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!\wrclk_control_slave_status_almostfull_q~q ),
	.datae(!\wrclk_control_slave_event_almostfull_q~q ),
	.dataf(!\wrclk_control_slave_ienable_register[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[2]~2 .extended_lut = "off";
defparam \wrclk_control_slave_read_mux[2]~2 .lut_mask = 64'h0040084804440C4C;
defparam \wrclk_control_slave_read_mux[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[2]~20 (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!\wrclk_control_slave_almostempty_threshold_register[2]~q ),
	.datad(!\wrclk_control_slave_read_mux[2]~2_combout ),
	.datae(!int_nxt_addr_reg_dly_2),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~1_sumout ),
	.datag(!\wrclk_control_slave_almostfull_threshold_register[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[2]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[2]~20 .extended_lut = "on";
defparam \wrclk_control_slave_read_mux[2]~20 .lut_mask = 64'h20FF02FFB9FF13FF;
defparam \wrclk_control_slave_read_mux[2]~20 .shared_arith = "off";

dffeas \wrclk_control_slave_almostempty_threshold_register[3] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_threshold_writedata[3]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\wrclk_control_slave_almostempty_threshold_register[3]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostempty_threshold_register[3] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostempty_threshold_register[3] .power_up = "low";

cyclonev_lcell_comb \LessThan2~0 (
	.dataa(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~17_sumout ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~21_sumout ),
	.datac(!\wrclk_control_slave_almostempty_threshold_register[0]~q ),
	.datad(!\wrclk_control_slave_almostempty_threshold_register[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~0 .extended_lut = "off";
defparam \LessThan2~0 .lut_mask = 64'h3701370137013701;
defparam \LessThan2~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan2~2 (
	.dataa(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~1_sumout ),
	.datab(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~5_sumout ),
	.datac(!\wrclk_control_slave_almostempty_threshold_register[2]~q ),
	.datad(!\wrclk_control_slave_almostempty_threshold_register[3]~q ),
	.datae(!\LessThan2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~2 .extended_lut = "off";
defparam \LessThan2~2 .lut_mask = 64'h7310F7317310F731;
defparam \LessThan2~2 .shared_arith = "off";

dffeas \wrclk_control_slave_almostempty_threshold_register[6] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_threshold_writedata[6]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\wrclk_control_slave_almostempty_threshold_register[6]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostempty_threshold_register[6] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostempty_threshold_register[6] .power_up = "low";

dffeas \wrclk_control_slave_almostempty_threshold_register[4] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_threshold_writedata[4]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\wrclk_control_slave_almostempty_threshold_register[4]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostempty_threshold_register[4] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostempty_threshold_register[4] .power_up = "low";

cyclonev_lcell_comb \LessThan2~3 (
	.dataa(!op_21),
	.datab(!\wrclk_control_slave_almostempty_threshold_register[6]~q ),
	.datac(!\wrclk_control_slave_almostempty_threshold_register[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~3 .extended_lut = "off";
defparam \LessThan2~3 .lut_mask = 64'hD4D4D4D4D4D4D4D4;
defparam \LessThan2~3 .shared_arith = "off";

dffeas \wrclk_control_slave_almostempty_threshold_register[7] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_threshold_writedata[7]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\wrclk_control_slave_almostempty_threshold_register[7]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostempty_threshold_register[7] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostempty_threshold_register[7] .power_up = "low";

dffeas \wrclk_control_slave_almostempty_threshold_register[5] (
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_threshold_writedata[5]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\wrclk_control_slave_almostempty_threshold_register[5]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_almostempty_threshold_register[5] .is_wysiwyg = "true";
defparam \wrclk_control_slave_almostempty_threshold_register[5] .power_up = "low";

cyclonev_lcell_comb \LessThan2~4 (
	.dataa(!op_21),
	.datab(!op_22),
	.datac(!\wrclk_control_slave_almostempty_threshold_register[6]~q ),
	.datad(!\wrclk_control_slave_almostempty_threshold_register[7]~q ),
	.datae(!op_2),
	.dataf(!\wrclk_control_slave_almostempty_threshold_register[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~4 .extended_lut = "off";
defparam \LessThan2~4 .lut_mask = 64'h08CE08CE8CEF08CE;
defparam \LessThan2~4 .shared_arith = "off";

cyclonev_lcell_comb \LessThan2~5 (
	.dataa(!op_21),
	.datab(!op_22),
	.datac(!\wrclk_control_slave_almostempty_threshold_register[6]~q ),
	.datad(!\wrclk_control_slave_almostempty_threshold_register[7]~q ),
	.datae(!op_2),
	.dataf(!\wrclk_control_slave_almostempty_threshold_register[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~5 .extended_lut = "off";
defparam \LessThan2~5 .lut_mask = 64'h8CAF00008CAF8CAF;
defparam \LessThan2~5 .shared_arith = "off";

cyclonev_lcell_comb \LessThan2~1 (
	.dataa(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~9_sumout ),
	.datab(!\LessThan2~2_combout ),
	.datac(!\LessThan2~3_combout ),
	.datad(!\LessThan2~4_combout ),
	.datae(!\LessThan2~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~1 .extended_lut = "off";
defparam \LessThan2~1 .lut_mask = 64'hFF001700FF001700;
defparam \LessThan2~1 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_status_almostempty_q~0 (
	.dataa(!\LessThan2~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_status_almostempty_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_status_almostempty_q~0 .extended_lut = "off";
defparam \wrclk_control_slave_status_almostempty_q~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wrclk_control_slave_status_almostempty_q~0 .shared_arith = "off";

dffeas wrclk_control_slave_status_almostempty_q(
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_status_almostempty_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_status_almostempty_q~q ),
	.prn(vcc));
defparam wrclk_control_slave_status_almostempty_q.is_wysiwyg = "true";
defparam wrclk_control_slave_status_almostempty_q.power_up = "low";

dffeas wrclk_control_slave_almostempty_n_reg(
	.clk(outclk_wire_0),
	.d(\LessThan2~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_almostempty_n_reg~q ),
	.prn(vcc));
defparam wrclk_control_slave_almostempty_n_reg.is_wysiwyg = "true";
defparam wrclk_control_slave_almostempty_n_reg.power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_event_almostempty_q~0 (
	.dataa(!\wrclk_control_slave_event_almostempty_q~q ),
	.datab(!\always7~0_combout ),
	.datac(!wrclk_control_slave_writedata[3]),
	.datad(!\LessThan2~1_combout ),
	.datae(!\wrclk_control_slave_almostempty_n_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_event_almostempty_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_event_almostempty_q~0 .extended_lut = "off";
defparam \wrclk_control_slave_event_almostempty_q~0 .lut_mask = 64'h5454FC545454FC54;
defparam \wrclk_control_slave_event_almostempty_q~0 .shared_arith = "off";

dffeas wrclk_control_slave_event_almostempty_q(
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_event_almostempty_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_event_almostempty_q~q ),
	.prn(vcc));
defparam wrclk_control_slave_event_almostempty_q.is_wysiwyg = "true";
defparam wrclk_control_slave_event_almostempty_q.power_up = "low";

dffeas \wrclk_control_slave_ienable_register[3] (
	.clk(outclk_wire_0),
	.d(wrclk_control_slave_writedata[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\wrclk_control_slave_ienable_register[3]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_ienable_register[3] .is_wysiwyg = "true";
defparam \wrclk_control_slave_ienable_register[3] .power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[3]~3 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!\wrclk_control_slave_status_almostempty_q~q ),
	.datae(!\wrclk_control_slave_event_almostempty_q~q ),
	.dataf(!\wrclk_control_slave_ienable_register[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[3]~3 .extended_lut = "off";
defparam \wrclk_control_slave_read_mux[3]~3 .lut_mask = 64'h0040084804440C4C;
defparam \wrclk_control_slave_read_mux[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[3]~16 (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!\wrclk_control_slave_almostempty_threshold_register[3]~q ),
	.datad(!\wrclk_control_slave_read_mux[3]~3_combout ),
	.datae(!int_nxt_addr_reg_dly_2),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~5_sumout ),
	.datag(!\wrclk_control_slave_almostfull_threshold_register[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[3]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[3]~16 .extended_lut = "on";
defparam \wrclk_control_slave_read_mux[3]~16 .lut_mask = 64'h20FF02FFB9FF13FF;
defparam \wrclk_control_slave_read_mux[3]~16 .shared_arith = "off";

cyclonev_lcell_comb wrclk_control_slave_status_overflow_signal(
	.dataa(!\the_dcfifo|wrfull~7_combout ),
	.datab(!m0_write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_status_overflow_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam wrclk_control_slave_status_overflow_signal.extended_lut = "off";
defparam wrclk_control_slave_status_overflow_signal.lut_mask = 64'h1111111111111111;
defparam wrclk_control_slave_status_overflow_signal.shared_arith = "off";

dffeas wrclk_control_slave_status_overflow_q(
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_status_overflow_signal~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_status_overflow_q~q ),
	.prn(vcc));
defparam wrclk_control_slave_status_overflow_q.is_wysiwyg = "true";
defparam wrclk_control_slave_status_overflow_q.power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_event_overflow_q~0 (
	.dataa(!\wrclk_control_slave_event_overflow_q~q ),
	.datab(!\always7~0_combout ),
	.datac(!wrclk_control_slave_writedata[4]),
	.datad(!\wrclk_control_slave_status_overflow_signal~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_event_overflow_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_event_overflow_q~0 .extended_lut = "off";
defparam \wrclk_control_slave_event_overflow_q~0 .lut_mask = 64'h54FC54FC54FC54FC;
defparam \wrclk_control_slave_event_overflow_q~0 .shared_arith = "off";

dffeas wrclk_control_slave_event_overflow_q(
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_event_overflow_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_event_overflow_q~q ),
	.prn(vcc));
defparam wrclk_control_slave_event_overflow_q.is_wysiwyg = "true";
defparam wrclk_control_slave_event_overflow_q.power_up = "low";

dffeas \wrclk_control_slave_ienable_register[4] (
	.clk(outclk_wire_0),
	.d(wrclk_control_slave_writedata[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\wrclk_control_slave_ienable_register[4]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_ienable_register[4] .is_wysiwyg = "true";
defparam \wrclk_control_slave_ienable_register[4] .power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[4]~4 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!\wrclk_control_slave_status_overflow_q~q ),
	.datae(!\wrclk_control_slave_event_overflow_q~q ),
	.dataf(!\wrclk_control_slave_ienable_register[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[4]~4 .extended_lut = "off";
defparam \wrclk_control_slave_read_mux[4]~4 .lut_mask = 64'h0040084804440C4C;
defparam \wrclk_control_slave_read_mux[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[4]~12 (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!\wrclk_control_slave_almostempty_threshold_register[4]~q ),
	.datad(!\wrclk_control_slave_read_mux[4]~4_combout ),
	.datae(!int_nxt_addr_reg_dly_2),
	.dataf(!\the_dcfifo|dual_clock_fifo|auto_generated|op_2~9_sumout ),
	.datag(!\wrclk_control_slave_almostfull_threshold_register[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[4]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[4]~12 .extended_lut = "on";
defparam \wrclk_control_slave_read_mux[4]~12 .lut_mask = 64'h20FF02FFB9FF13FF;
defparam \wrclk_control_slave_read_mux[4]~12 .shared_arith = "off";

cyclonev_lcell_comb wrclk_control_slave_status_underflow_signal(
	.dataa(!\the_dcfifo|dual_clock_fifo|auto_generated|wrempty_eq_comp|aneb_result_wire[0]~combout ),
	.datab(!\rdreq_sync_i|dreg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_status_underflow_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam wrclk_control_slave_status_underflow_signal.extended_lut = "off";
defparam wrclk_control_slave_status_underflow_signal.lut_mask = 64'h2222222222222222;
defparam wrclk_control_slave_status_underflow_signal.shared_arith = "off";

dffeas wrclk_control_slave_status_underflow_q(
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_status_underflow_signal~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_status_underflow_q~q ),
	.prn(vcc));
defparam wrclk_control_slave_status_underflow_q.is_wysiwyg = "true";
defparam wrclk_control_slave_status_underflow_q.power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_event_underflow_q~0 (
	.dataa(!\wrclk_control_slave_event_underflow_q~q ),
	.datab(!\always7~0_combout ),
	.datac(!wrclk_control_slave_writedata[5]),
	.datad(!\wrclk_control_slave_status_underflow_signal~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_event_underflow_q~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_event_underflow_q~0 .extended_lut = "off";
defparam \wrclk_control_slave_event_underflow_q~0 .lut_mask = 64'h54FC54FC54FC54FC;
defparam \wrclk_control_slave_event_underflow_q~0 .shared_arith = "off";

dffeas wrclk_control_slave_event_underflow_q(
	.clk(outclk_wire_0),
	.d(\wrclk_control_slave_event_underflow_q~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wrclk_control_slave_event_underflow_q~q ),
	.prn(vcc));
defparam wrclk_control_slave_event_underflow_q.is_wysiwyg = "true";
defparam wrclk_control_slave_event_underflow_q.power_up = "low";

dffeas \wrclk_control_slave_ienable_register[5] (
	.clk(outclk_wire_0),
	.d(wrclk_control_slave_writedata[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\wrclk_control_slave_ienable_register[5]~q ),
	.prn(vcc));
defparam \wrclk_control_slave_ienable_register[5] .is_wysiwyg = "true";
defparam \wrclk_control_slave_ienable_register[5] .power_up = "low";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[5]~5 (
	.dataa(!int_nxt_addr_reg_dly_2),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(!\wrclk_control_slave_status_underflow_q~q ),
	.datae(!\wrclk_control_slave_event_underflow_q~q ),
	.dataf(!\wrclk_control_slave_ienable_register[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[5]~5 .extended_lut = "off";
defparam \wrclk_control_slave_read_mux[5]~5 .lut_mask = 64'h0040084804440C4C;
defparam \wrclk_control_slave_read_mux[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[5]~8 (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_4),
	.datac(!\wrclk_control_slave_almostempty_threshold_register[5]~q ),
	.datad(!\wrclk_control_slave_read_mux[5]~5_combout ),
	.datae(!int_nxt_addr_reg_dly_2),
	.dataf(!op_2),
	.datag(!\wrclk_control_slave_almostfull_threshold_register[5]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[5]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[5]~8 .extended_lut = "on";
defparam \wrclk_control_slave_read_mux[5]~8 .lut_mask = 64'h20FF02FFB9FF13FF;
defparam \wrclk_control_slave_read_mux[5]~8 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[6]~6 (
	.dataa(!op_21),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\wrclk_control_slave_almostfull_threshold_register[6]~q ),
	.dataf(!\wrclk_control_slave_almostempty_threshold_register[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[6]~6 .extended_lut = "off";
defparam \wrclk_control_slave_read_mux[6]~6 .lut_mask = 64'h4C0540054F054305;
defparam \wrclk_control_slave_read_mux[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \wrclk_control_slave_read_mux[7]~7 (
	.dataa(!op_22),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!int_nxt_addr_reg_dly_4),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!\wrclk_control_slave_almostfull_threshold_register[7]~q ),
	.dataf(!\wrclk_control_slave_almostempty_threshold_register[7]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrclk_control_slave_read_mux[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrclk_control_slave_read_mux[7]~7 .extended_lut = "off";
defparam \wrclk_control_slave_read_mux[7]~7 .lut_mask = 64'h4C0540054F054305;
defparam \wrclk_control_slave_read_mux[7]~7 .shared_arith = "off";

endmodule

module Computer_System_altera_std_synchronizer (
	clk,
	reset_n,
	dreg_2,
	din)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	reset_n;
output 	dreg_2;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;
wire \dreg[1]~q ;


dffeas \dreg[2] (
	.clk(clk),
	.d(\dreg[1]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_2),
	.prn(vcc));
defparam \dreg[2] .is_wysiwyg = "true";
defparam \dreg[2] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[1]~q ),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

endmodule

module Computer_System_altera_std_synchronizer_1 (
	din,
	reset_n,
	dreg_2,
	clk)/* synthesis synthesis_greybox=0 */;
input 	din;
input 	reset_n;
output 	dreg_2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;
wire \dreg[1]~q ;


dffeas \dreg[2] (
	.clk(clk),
	.d(\dreg[1]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_2),
	.prn(vcc));
defparam \dreg[2] .is_wysiwyg = "true";
defparam \dreg[2] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[1]~q ),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

endmodule

module Computer_System_Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	outclk_wire_0,
	op_2,
	op_21,
	op_22,
	op_23,
	op_24,
	op_25,
	op_26,
	op_27,
	op_1,
	op_11,
	op_12,
	op_13,
	op_14,
	op_15,
	op_16,
	op_17,
	data_wire_2,
	aneb_result_wire_0,
	aneb_result_wire_01,
	aneb_result_wire_02,
	aneb_result_wire_03,
	wrfull,
	wrfull1,
	wrfull2,
	m0_write,
	in_data_reg_0,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	wrfull3,
	wrfull4,
	comb,
	aneb_result_wire_04,
	rdfull,
	rdfull1,
	rdfull2,
	wrfull5,
	aneb_result_wire_05,
	fifo_hps_to_fpga_out_read,
	clock_bridge_0_in_clk_clk)/* synthesis synthesis_greybox=0 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
input 	outclk_wire_0;
output 	op_2;
output 	op_21;
output 	op_22;
output 	op_23;
output 	op_24;
output 	op_25;
output 	op_26;
output 	op_27;
output 	op_1;
output 	op_11;
output 	op_12;
output 	op_13;
output 	op_14;
output 	op_15;
output 	op_16;
output 	op_17;
output 	data_wire_2;
output 	aneb_result_wire_0;
output 	aneb_result_wire_01;
output 	aneb_result_wire_02;
output 	aneb_result_wire_03;
output 	wrfull;
output 	wrfull1;
output 	wrfull2;
input 	m0_write;
input 	in_data_reg_0;
input 	in_data_reg_1;
input 	in_data_reg_2;
input 	in_data_reg_3;
input 	in_data_reg_4;
input 	in_data_reg_5;
input 	in_data_reg_6;
input 	in_data_reg_7;
input 	in_data_reg_8;
input 	in_data_reg_9;
input 	in_data_reg_10;
input 	in_data_reg_11;
input 	in_data_reg_12;
input 	in_data_reg_13;
input 	in_data_reg_14;
input 	in_data_reg_15;
input 	in_data_reg_16;
input 	in_data_reg_17;
input 	in_data_reg_18;
input 	in_data_reg_19;
input 	in_data_reg_20;
input 	in_data_reg_21;
input 	in_data_reg_22;
input 	in_data_reg_23;
input 	in_data_reg_24;
input 	in_data_reg_25;
input 	in_data_reg_26;
input 	in_data_reg_27;
input 	in_data_reg_28;
input 	in_data_reg_29;
input 	in_data_reg_30;
input 	in_data_reg_31;
output 	wrfull3;
output 	wrfull4;
input 	comb;
output 	aneb_result_wire_04;
output 	rdfull;
output 	rdfull1;
output 	rdfull2;
output 	wrfull5;
output 	aneb_result_wire_05;
input 	fifo_hps_to_fpga_out_read;
input 	clock_bridge_0_in_clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dual_clock_fifo|auto_generated|wraclr|dffe13a[0]~q ;
wire \dual_clock_fifo|auto_generated|wrptr_g[1]~q ;
wire \dual_clock_fifo|auto_generated|ws_dgrp|dffpipe18|dffe20a[1]~q ;
wire \dual_clock_fifo|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~0_combout ;
wire \dual_clock_fifo|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~1_combout ;
wire \dual_clock_fifo|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~2_combout ;
wire \wrfull~3_combout ;
wire \wrfull~6_combout ;


Computer_System_dcfifo_1 dual_clock_fifo(
	.q({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wrclk(outclk_wire_0),
	.op_2(op_2),
	.op_21(op_21),
	.op_22(op_22),
	.op_23(op_23),
	.op_24(op_24),
	.op_25(op_25),
	.op_26(op_26),
	.op_27(op_27),
	.op_1(op_1),
	.op_11(op_11),
	.op_12(op_12),
	.op_13(op_13),
	.op_14(op_14),
	.op_15(op_15),
	.op_16(op_16),
	.op_17(op_17),
	.data_wire_2(data_wire_2),
	.aneb_result_wire_0(aneb_result_wire_0),
	.aneb_result_wire_01(aneb_result_wire_01),
	.aneb_result_wire_02(aneb_result_wire_02),
	.aneb_result_wire_03(aneb_result_wire_03),
	.wrfull(wrfull),
	.wrfull1(wrfull1),
	.dffe13a_0(\dual_clock_fifo|auto_generated|wraclr|dffe13a[0]~q ),
	.wrptr_g_1(\dual_clock_fifo|auto_generated|wrptr_g[1]~q ),
	.dffe20a_1(\dual_clock_fifo|auto_generated|ws_dgrp|dffpipe18|dffe20a[1]~q ),
	.aneb_result_wire_04(\dual_clock_fifo|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~0_combout ),
	.aneb_result_wire_05(\dual_clock_fifo|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~1_combout ),
	.aneb_result_wire_06(\dual_clock_fifo|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~2_combout ),
	.wrfull2(wrfull2),
	.m0_write(m0_write),
	.data({in_data_reg_31,in_data_reg_30,in_data_reg_29,in_data_reg_28,in_data_reg_27,in_data_reg_26,in_data_reg_25,in_data_reg_24,in_data_reg_23,in_data_reg_22,in_data_reg_21,in_data_reg_20,in_data_reg_19,in_data_reg_18,in_data_reg_17,in_data_reg_16,in_data_reg_15,in_data_reg_14,
in_data_reg_13,in_data_reg_12,in_data_reg_11,in_data_reg_10,in_data_reg_9,in_data_reg_8,in_data_reg_7,in_data_reg_6,in_data_reg_5,in_data_reg_4,in_data_reg_3,in_data_reg_2,in_data_reg_1,in_data_reg_0}),
	.wrfull3(wrfull4),
	.comb(comb),
	.aneb_result_wire_07(aneb_result_wire_04),
	.aneb_result_wire_08(aneb_result_wire_05),
	.fifo_hps_to_fpga_out_read(fifo_hps_to_fpga_out_read),
	.rdclk(clock_bridge_0_in_clk_clk));

cyclonev_lcell_comb \wrfull~0 (
	.dataa(!op_2),
	.datab(!op_21),
	.datac(!op_22),
	.datad(!op_23),
	.datae(!op_24),
	.dataf(!op_25),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wrfull),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrfull~0 .extended_lut = "off";
defparam \wrfull~0 .lut_mask = 64'h0000000100010001;
defparam \wrfull~0 .shared_arith = "off";

cyclonev_lcell_comb \wrfull~1 (
	.dataa(!op_26),
	.datab(!op_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wrfull1),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrfull~1 .extended_lut = "off";
defparam \wrfull~1 .lut_mask = 64'h1111111111111111;
defparam \wrfull~1 .shared_arith = "off";

cyclonev_lcell_comb \wrfull~2 (
	.dataa(!\dual_clock_fifo|auto_generated|wraclr|dffe13a[0]~q ),
	.datab(!\dual_clock_fifo|auto_generated|wrptr_g[1]~q ),
	.datac(!\dual_clock_fifo|auto_generated|ws_dgrp|dffpipe18|dffe20a[1]~q ),
	.datad(!\dual_clock_fifo|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~0_combout ),
	.datae(!\dual_clock_fifo|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~1_combout ),
	.dataf(!\dual_clock_fifo|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wrfull2),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrfull~2 .extended_lut = "off";
defparam \wrfull~2 .lut_mask = 64'h5555555555555514;
defparam \wrfull~2 .shared_arith = "off";

cyclonev_lcell_comb \wrfull~4 (
	.dataa(!op_21),
	.datab(!op_22),
	.datac(!op_23),
	.datad(!op_26),
	.datae(!op_27),
	.dataf(!\wrfull~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wrfull3),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrfull~4 .extended_lut = "off";
defparam \wrfull~4 .lut_mask = 64'h0000000000000001;
defparam \wrfull~4 .shared_arith = "off";

cyclonev_lcell_comb \wrfull~5 (
	.dataa(!op_2),
	.datab(!op_21),
	.datac(!op_22),
	.datad(!op_24),
	.datae(!op_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wrfull4),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrfull~5 .extended_lut = "off";
defparam \wrfull~5 .lut_mask = 64'h0001010100010101;
defparam \wrfull~5 .shared_arith = "off";

cyclonev_lcell_comb \rdfull~0 (
	.dataa(!op_1),
	.datab(!op_11),
	.datac(!op_12),
	.datad(!op_13),
	.datae(!op_14),
	.dataf(!op_15),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rdfull),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdfull~0 .extended_lut = "off";
defparam \rdfull~0 .lut_mask = 64'h0000000000000007;
defparam \rdfull~0 .shared_arith = "off";

cyclonev_lcell_comb \rdfull~1 (
	.dataa(!op_16),
	.datab(!op_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rdfull1),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdfull~1 .extended_lut = "off";
defparam \rdfull~1 .lut_mask = 64'h1111111111111111;
defparam \rdfull~1 .shared_arith = "off";

cyclonev_lcell_comb \rdfull~2 (
	.dataa(!aneb_result_wire_04),
	.datab(!rdfull),
	.datac(!rdfull1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rdfull2),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdfull~2 .extended_lut = "off";
defparam \rdfull~2 .lut_mask = 64'h5757575757575757;
defparam \rdfull~2 .shared_arith = "off";

cyclonev_lcell_comb \wrfull~7 (
	.dataa(!op_22),
	.datab(!op_23),
	.datac(!op_26),
	.datad(!op_27),
	.datae(!\wrfull~6_combout ),
	.dataf(!wrfull2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wrfull5),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrfull~7 .extended_lut = "off";
defparam \wrfull~7 .lut_mask = 64'hFFFFFFFF00000001;
defparam \wrfull~7 .shared_arith = "off";

cyclonev_lcell_comb \wrfull~3 (
	.dataa(!op_2),
	.datab(!op_24),
	.datac(!op_25),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrfull~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrfull~3 .extended_lut = "off";
defparam \wrfull~3 .lut_mask = 64'h1515151515151515;
defparam \wrfull~3 .shared_arith = "off";

cyclonev_lcell_comb \wrfull~6 (
	.dataa(!op_2),
	.datab(!op_21),
	.datac(!op_24),
	.datad(!op_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrfull~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrfull~6 .extended_lut = "off";
defparam \wrfull~6 .lut_mask = 64'h0111011101110111;
defparam \wrfull~6 .shared_arith = "off";

endmodule

module Computer_System_dcfifo_1 (
	q,
	wrclk,
	op_2,
	op_21,
	op_22,
	op_23,
	op_24,
	op_25,
	op_26,
	op_27,
	op_1,
	op_11,
	op_12,
	op_13,
	op_14,
	op_15,
	op_16,
	op_17,
	data_wire_2,
	aneb_result_wire_0,
	aneb_result_wire_01,
	aneb_result_wire_02,
	aneb_result_wire_03,
	wrfull,
	wrfull1,
	dffe13a_0,
	wrptr_g_1,
	dffe20a_1,
	aneb_result_wire_04,
	aneb_result_wire_05,
	aneb_result_wire_06,
	wrfull2,
	m0_write,
	data,
	wrfull3,
	comb,
	aneb_result_wire_07,
	aneb_result_wire_08,
	fifo_hps_to_fpga_out_read,
	rdclk)/* synthesis synthesis_greybox=0 */;
output 	[31:0] q;
input 	wrclk;
output 	op_2;
output 	op_21;
output 	op_22;
output 	op_23;
output 	op_24;
output 	op_25;
output 	op_26;
output 	op_27;
output 	op_1;
output 	op_11;
output 	op_12;
output 	op_13;
output 	op_14;
output 	op_15;
output 	op_16;
output 	op_17;
output 	data_wire_2;
output 	aneb_result_wire_0;
output 	aneb_result_wire_01;
output 	aneb_result_wire_02;
output 	aneb_result_wire_03;
input 	wrfull;
input 	wrfull1;
output 	dffe13a_0;
output 	wrptr_g_1;
output 	dffe20a_1;
output 	aneb_result_wire_04;
output 	aneb_result_wire_05;
output 	aneb_result_wire_06;
input 	wrfull2;
input 	m0_write;
input 	[31:0] data;
input 	wrfull3;
input 	comb;
output 	aneb_result_wire_07;
output 	aneb_result_wire_08;
input 	fifo_hps_to_fpga_out_read;
input 	rdclk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_dcfifo_k482 auto_generated(
	.q({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.wrclk(wrclk),
	.op_2(op_2),
	.op_21(op_21),
	.op_22(op_22),
	.op_23(op_23),
	.op_24(op_24),
	.op_25(op_25),
	.op_26(op_26),
	.op_27(op_27),
	.op_1(op_1),
	.op_11(op_11),
	.op_12(op_12),
	.op_13(op_13),
	.op_14(op_14),
	.op_15(op_15),
	.op_16(op_16),
	.op_17(op_17),
	.data_wire_2(data_wire_2),
	.aneb_result_wire_0(aneb_result_wire_0),
	.aneb_result_wire_01(aneb_result_wire_01),
	.aneb_result_wire_02(aneb_result_wire_02),
	.aneb_result_wire_03(aneb_result_wire_03),
	.wrfull(wrfull),
	.wrfull1(wrfull1),
	.dffe13a_0(dffe13a_0),
	.wrptr_g_1(wrptr_g_1),
	.dffe20a_1(dffe20a_1),
	.aneb_result_wire_04(aneb_result_wire_04),
	.aneb_result_wire_05(aneb_result_wire_05),
	.aneb_result_wire_06(aneb_result_wire_06),
	.wrfull2(wrfull2),
	.m0_write(m0_write),
	.data({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.wrfull3(wrfull3),
	.comb(comb),
	.aneb_result_wire_07(aneb_result_wire_07),
	.aneb_result_wire_08(aneb_result_wire_08),
	.fifo_hps_to_fpga_out_read(fifo_hps_to_fpga_out_read),
	.rdclk(rdclk));

endmodule

module Computer_System_dcfifo_k482 (
	q,
	wrclk,
	op_2,
	op_21,
	op_22,
	op_23,
	op_24,
	op_25,
	op_26,
	op_27,
	op_1,
	op_11,
	op_12,
	op_13,
	op_14,
	op_15,
	op_16,
	op_17,
	data_wire_2,
	aneb_result_wire_0,
	aneb_result_wire_01,
	aneb_result_wire_02,
	aneb_result_wire_03,
	wrfull,
	wrfull1,
	dffe13a_0,
	wrptr_g_1,
	dffe20a_1,
	aneb_result_wire_04,
	aneb_result_wire_05,
	aneb_result_wire_06,
	wrfull2,
	m0_write,
	data,
	wrfull3,
	comb,
	aneb_result_wire_07,
	aneb_result_wire_08,
	fifo_hps_to_fpga_out_read,
	rdclk)/* synthesis synthesis_greybox=0 */;
output 	[31:0] q;
input 	wrclk;
output 	op_2;
output 	op_21;
output 	op_22;
output 	op_23;
output 	op_24;
output 	op_25;
output 	op_26;
output 	op_27;
output 	op_1;
output 	op_11;
output 	op_12;
output 	op_13;
output 	op_14;
output 	op_15;
output 	op_16;
output 	op_17;
output 	data_wire_2;
output 	aneb_result_wire_0;
output 	aneb_result_wire_01;
output 	aneb_result_wire_02;
output 	aneb_result_wire_03;
input 	wrfull;
input 	wrfull1;
output 	dffe13a_0;
output 	wrptr_g_1;
output 	dffe20a_1;
output 	aneb_result_wire_04;
output 	aneb_result_wire_05;
output 	aneb_result_wire_06;
input 	wrfull2;
input 	m0_write;
input 	[31:0] data;
input 	wrfull3;
input 	comb;
output 	aneb_result_wire_07;
output 	aneb_result_wire_08;
input 	fifo_hps_to_fpga_out_read;
input 	rdclk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \rdptr_g[1]~q ;
wire \rs_dgwp|dffpipe15|dffe17a[1]~q ;
wire \rdptr_g[6]~q ;
wire \rs_dgwp|dffpipe15|dffe17a[6]~q ;
wire \rdptr_g[4]~q ;
wire \rs_dgwp|dffpipe15|dffe17a[4]~q ;
wire \rdptr_g[5]~q ;
wire \rs_dgwp|dffpipe15|dffe17a[5]~q ;
wire \rdptr_g[2]~q ;
wire \rs_dgwp|dffpipe15|dffe17a[2]~q ;
wire \rdptr_g[3]~q ;
wire \rs_dgwp|dffpipe15|dffe17a[3]~q ;
wire \rdptr_g[0]~q ;
wire \rs_dgwp|dffpipe15|dffe17a[0]~q ;
wire \rdptr_g[8]~q ;
wire \rs_dgwp|dffpipe15|dffe17a[8]~q ;
wire \rdptr_g[7]~q ;
wire \rs_dgwp|dffpipe15|dffe17a[7]~q ;
wire \wrptr_g[6]~q ;
wire \ws_dgrp|dffpipe18|dffe20a[6]~q ;
wire \wrptr_g[4]~q ;
wire \ws_dgrp|dffpipe18|dffe20a[4]~q ;
wire \wrptr_g[5]~q ;
wire \ws_dgrp|dffpipe18|dffe20a[5]~q ;
wire \wrptr_g[2]~q ;
wire \ws_dgrp|dffpipe18|dffe20a[2]~q ;
wire \wrptr_g[3]~q ;
wire \ws_dgrp|dffpipe18|dffe20a[3]~q ;
wire \wrptr_g[0]~q ;
wire \ws_dgrp|dffpipe18|dffe20a[0]~q ;
wire \wrptr_g[8]~q ;
wire \ws_dgrp|dffpipe18|dffe20a[8]~q ;
wire \wrptr_g[7]~q ;
wire \ws_dgrp|dffpipe18|dffe20a[7]~q ;
wire \wrptr_g1p|_~0_combout ;
wire \rdaclr|dffe13a[0]~q ;
wire \valid_rdreq~0_combout ;
wire \ram_address_a[7]~combout ;
wire \rdptr_g1p|counter5a0~q ;
wire \rdptr_g1p|counter5a1~q ;
wire \rdptr_g1p|counter5a2~q ;
wire \rdptr_g1p|counter5a3~q ;
wire \rdptr_g1p|counter5a4~q ;
wire \rdptr_g1p|counter5a5~q ;
wire \rdptr_g1p|counter5a6~q ;
wire \rdptr_g1p|counter5a7~q ;
wire \rdptr_g1p|counter5a8~q ;
wire \rdptr_g1p|_~0_combout ;
wire \ws_brp|dffe14a[2]~q ;
wire \ws_bwp|dffe14a[2]~q ;
wire \ws_brp|dffe14a[3]~q ;
wire \ws_bwp|dffe14a[3]~q ;
wire \ws_brp|dffe14a[4]~q ;
wire \ws_bwp|dffe14a[4]~q ;
wire \ws_brp|dffe14a[5]~q ;
wire \ws_bwp|dffe14a[5]~q ;
wire \ws_brp|dffe14a[0]~q ;
wire \ws_bwp|dffe14a[0]~q ;
wire \ws_brp|dffe14a[1]~q ;
wire \ws_bwp|dffe14a[1]~q ;
wire \ws_brp|dffe14a[6]~q ;
wire \ws_bwp|dffe14a[6]~q ;
wire \ws_brp|dffe14a[7]~q ;
wire \ws_bwp|dffe14a[7]~q ;
wire \wrptr_g1p|counter8a1~q ;
wire \wrptr_g1p|counter8a6~q ;
wire \wrptr_g1p|counter8a4~q ;
wire \wrptr_g1p|counter8a5~q ;
wire \wrptr_g1p|counter8a2~q ;
wire \wrptr_g1p|counter8a3~q ;
wire \wrptr_g1p|counter8a0~q ;
wire \wrptr_g1p|counter8a8~q ;
wire \wrptr_g1p|counter8a7~q ;
wire \delayed_wrptr_g[1]~q ;
wire \delayed_wrptr_g[6]~q ;
wire \delayed_wrptr_g[4]~q ;
wire \delayed_wrptr_g[5]~q ;
wire \delayed_wrptr_g[2]~q ;
wire \delayed_wrptr_g[3]~q ;
wire \delayed_wrptr_g[0]~q ;
wire \delayed_wrptr_g[8]~q ;
wire \delayed_wrptr_g[7]~q ;
wire \rs_brp|dffe14a[0]~q ;
wire \rs_bwp|dffe14a[0]~q ;
wire \rs_brp|dffe14a[1]~q ;
wire \rs_bwp|dffe14a[1]~q ;
wire \rs_brp|dffe14a[2]~q ;
wire \rs_bwp|dffe14a[2]~q ;
wire \rs_brp|dffe14a[3]~q ;
wire \rs_bwp|dffe14a[3]~q ;
wire \rs_brp|dffe14a[4]~q ;
wire \rs_bwp|dffe14a[4]~q ;
wire \rs_brp|dffe14a[5]~q ;
wire \rs_bwp|dffe14a[5]~q ;
wire \rs_brp|dffe14a[6]~q ;
wire \rs_bwp|dffe14a[6]~q ;
wire \rs_brp|dffe14a[7]~q ;
wire \rs_bwp|dffe14a[7]~q ;
wire \ws_dgrp_gray2bin|xor7~combout ;
wire \ws_dgrp_gray2bin|xor6~combout ;
wire \ws_dgrp_gray2bin|xor5~combout ;
wire \ws_dgrp_gray2bin|xor4~combout ;
wire \ws_dgrp_gray2bin|xor3~combout ;
wire \ws_dgrp_gray2bin|xor2~combout ;
wire \wrptr_g_gray2bin|xor6~combout ;
wire \wrptr_g_gray2bin|xor5~combout ;
wire \wrptr_g_gray2bin|xor4~combout ;
wire \wrptr_g_gray2bin|xor3~combout ;
wire \wrptr_g_gray2bin|xor2~combout ;
wire \ws_dgrp_gray2bin|xor1~combout ;
wire \ws_dgrp_gray2bin|xor0~combout ;
wire \wrptr_g_gray2bin|xor1~combout ;
wire \wrptr_g_gray2bin|xor0~combout ;
wire \rdptr_g_gray2bin|xor7~combout ;
wire \rdptr_g_gray2bin|xor3~combout ;
wire \rdptr_g_gray2bin|xor0~combout ;
wire \rs_dgwp_gray2bin|xor7~combout ;
wire \rs_dgwp_gray2bin|xor3~combout ;
wire \rs_dgwp_gray2bin|xor0~combout ;
wire \rdptr_g_gray2bin|xor1~combout ;
wire \rs_dgwp_gray2bin|xor1~combout ;
wire \rdptr_g_gray2bin|xor2~combout ;
wire \rs_dgwp_gray2bin|xor2~combout ;
wire \rdptr_g_gray2bin|xor6~combout ;
wire \rdptr_g_gray2bin|xor4~combout ;
wire \rs_dgwp_gray2bin|xor6~combout ;
wire \rs_dgwp_gray2bin|xor4~combout ;
wire \rdptr_g_gray2bin|xor5~combout ;
wire \rs_dgwp_gray2bin|xor5~combout ;
wire \rdptr_g[0]~0_combout ;
wire \wrptr_g[0]~0_combout ;
wire \rdptr_g1p|counter5a0~_wirecell_combout ;
wire \op_2~2 ;
wire \op_2~3 ;
wire \op_2~6 ;
wire \op_2~7 ;
wire \op_2~10 ;
wire \op_2~11 ;
wire \op_2~14 ;
wire \op_2~15 ;
wire \op_2~18 ;
wire \op_2~19 ;
wire \op_2~22 ;
wire \op_2~23 ;
wire \op_2~26 ;
wire \op_2~27 ;
wire \op_1~2 ;
wire \op_1~3 ;
wire \op_1~6 ;
wire \op_1~7 ;
wire \op_1~10 ;
wire \op_1~11 ;
wire \op_1~14 ;
wire \op_1~15 ;
wire \op_1~18 ;
wire \op_1~19 ;
wire \op_1~22 ;
wire \op_1~23 ;
wire \op_1~26 ;
wire \op_1~27 ;


Computer_System_cmpr_1v5_3 wrfull_eq_comp(
	.wrptr_g_6(\wrptr_g[6]~q ),
	.dffe20a_6(\ws_dgrp|dffpipe18|dffe20a[6]~q ),
	.wrptr_g_4(\wrptr_g[4]~q ),
	.dffe20a_4(\ws_dgrp|dffpipe18|dffe20a[4]~q ),
	.wrptr_g_5(\wrptr_g[5]~q ),
	.dffe20a_5(\ws_dgrp|dffpipe18|dffe20a[5]~q ),
	.aneb_result_wire_0(aneb_result_wire_04),
	.wrptr_g_2(\wrptr_g[2]~q ),
	.dffe20a_2(\ws_dgrp|dffpipe18|dffe20a[2]~q ),
	.wrptr_g_3(\wrptr_g[3]~q ),
	.dffe20a_3(\ws_dgrp|dffpipe18|dffe20a[3]~q ),
	.wrptr_g_0(\wrptr_g[0]~q ),
	.dffe20a_0(\ws_dgrp|dffpipe18|dffe20a[0]~q ),
	.aneb_result_wire_01(aneb_result_wire_05),
	.wrptr_g_8(\wrptr_g[8]~q ),
	.dffe20a_8(\ws_dgrp|dffpipe18|dffe20a[8]~q ),
	.wrptr_g_7(\wrptr_g[7]~q ),
	.dffe20a_7(\ws_dgrp|dffpipe18|dffe20a[7]~q ),
	.aneb_result_wire_02(aneb_result_wire_06));

Computer_System_cmpr_1v5_2 wrempty_eq_comp(
	.wrptr_g_1(wrptr_g_1),
	.dffe20a_1(dffe20a_1),
	.aneb_result_wire_0(aneb_result_wire_04),
	.aneb_result_wire_01(aneb_result_wire_05),
	.wrptr_g_8(\wrptr_g[8]~q ),
	.dffe20a_8(\ws_dgrp|dffpipe18|dffe20a[8]~q ),
	.wrptr_g_7(\wrptr_g[7]~q ),
	.dffe20a_7(\ws_dgrp|dffpipe18|dffe20a[7]~q ),
	.aneb_result_wire_02(aneb_result_wire_08));

Computer_System_cmpr_1v5_1 rdfull_eq_comp(
	.data_wire_2(data_wire_2),
	.rdptr_g_6(\rdptr_g[6]~q ),
	.dffe17a_6(\rs_dgwp|dffpipe15|dffe17a[6]~q ),
	.rdptr_g_4(\rdptr_g[4]~q ),
	.dffe17a_4(\rs_dgwp|dffpipe15|dffe17a[4]~q ),
	.rdptr_g_5(\rdptr_g[5]~q ),
	.dffe17a_5(\rs_dgwp|dffpipe15|dffe17a[5]~q ),
	.aneb_result_wire_0(aneb_result_wire_0),
	.rdptr_g_2(\rdptr_g[2]~q ),
	.dffe17a_2(\rs_dgwp|dffpipe15|dffe17a[2]~q ),
	.rdptr_g_3(\rdptr_g[3]~q ),
	.dffe17a_3(\rs_dgwp|dffpipe15|dffe17a[3]~q ),
	.rdptr_g_0(\rdptr_g[0]~q ),
	.dffe17a_0(\rs_dgwp|dffpipe15|dffe17a[0]~q ),
	.aneb_result_wire_01(aneb_result_wire_01),
	.rdptr_g_8(\rdptr_g[8]~q ),
	.dffe17a_8(\rs_dgwp|dffpipe15|dffe17a[8]~q ),
	.rdptr_g_7(\rdptr_g[7]~q ),
	.dffe17a_7(\rs_dgwp|dffpipe15|dffe17a[7]~q ),
	.aneb_result_wire_02(aneb_result_wire_07));

Computer_System_cmpr_1v5 rdempty_eq_comp(
	.rdptr_g_1(\rdptr_g[1]~q ),
	.dffe17a_1(\rs_dgwp|dffpipe15|dffe17a[1]~q ),
	.data_wire_2(data_wire_2),
	.aneb_result_wire_0(aneb_result_wire_0),
	.aneb_result_wire_01(aneb_result_wire_01),
	.rdptr_g_8(\rdptr_g[8]~q ),
	.dffe17a_8(\rs_dgwp|dffpipe15|dffe17a[8]~q ),
	.rdptr_g_7(\rdptr_g[7]~q ),
	.dffe17a_7(\rs_dgwp|dffpipe15|dffe17a[7]~q ),
	.aneb_result_wire_02(aneb_result_wire_02),
	.aneb_result_wire_03(aneb_result_wire_03));

Computer_System_alt_synch_pipe_1ol ws_dgrp(
	.clock(wrclk),
	.rdptr_g_1(\rdptr_g[1]~q ),
	.rdptr_g_6(\rdptr_g[6]~q ),
	.rdptr_g_4(\rdptr_g[4]~q ),
	.rdptr_g_5(\rdptr_g[5]~q ),
	.rdptr_g_2(\rdptr_g[2]~q ),
	.rdptr_g_3(\rdptr_g[3]~q ),
	.rdptr_g_0(\rdptr_g[0]~q ),
	.rdptr_g_8(\rdptr_g[8]~q ),
	.rdptr_g_7(\rdptr_g[7]~q ),
	.clrn(dffe13a_0),
	.dffe20a_1(dffe20a_1),
	.dffe20a_6(\ws_dgrp|dffpipe18|dffe20a[6]~q ),
	.dffe20a_4(\ws_dgrp|dffpipe18|dffe20a[4]~q ),
	.dffe20a_5(\ws_dgrp|dffpipe18|dffe20a[5]~q ),
	.dffe20a_2(\ws_dgrp|dffpipe18|dffe20a[2]~q ),
	.dffe20a_3(\ws_dgrp|dffpipe18|dffe20a[3]~q ),
	.dffe20a_0(\ws_dgrp|dffpipe18|dffe20a[0]~q ),
	.dffe20a_8(\ws_dgrp|dffpipe18|dffe20a[8]~q ),
	.dffe20a_7(\ws_dgrp|dffpipe18|dffe20a[7]~q ));

Computer_System_dffpipe_gd9_3 ws_bwp(
	.clock(wrclk),
	.clrn(dffe13a_0),
	.ram_address_a_7(\ram_address_a[7]~combout ),
	.dffe14a_2(\ws_bwp|dffe14a[2]~q ),
	.dffe14a_3(\ws_bwp|dffe14a[3]~q ),
	.dffe14a_4(\ws_bwp|dffe14a[4]~q ),
	.dffe14a_5(\ws_bwp|dffe14a[5]~q ),
	.dffe14a_0(\ws_bwp|dffe14a[0]~q ),
	.dffe14a_1(\ws_bwp|dffe14a[1]~q ),
	.dffe14a_6(\ws_bwp|dffe14a[6]~q ),
	.dffe14a_7(\ws_bwp|dffe14a[7]~q ),
	.xor6(\wrptr_g_gray2bin|xor6~combout ),
	.xor5(\wrptr_g_gray2bin|xor5~combout ),
	.xor4(\wrptr_g_gray2bin|xor4~combout ),
	.xor3(\wrptr_g_gray2bin|xor3~combout ),
	.xor2(\wrptr_g_gray2bin|xor2~combout ),
	.xor1(\wrptr_g_gray2bin|xor1~combout ),
	.xor0(\wrptr_g_gray2bin|xor0~combout ));

Computer_System_dffpipe_gd9_2 ws_brp(
	.clock(wrclk),
	.clrn(dffe13a_0),
	.dffe14a_2(\ws_brp|dffe14a[2]~q ),
	.dffe14a_3(\ws_brp|dffe14a[3]~q ),
	.dffe14a_4(\ws_brp|dffe14a[4]~q ),
	.dffe14a_5(\ws_brp|dffe14a[5]~q ),
	.dffe14a_0(\ws_brp|dffe14a[0]~q ),
	.dffe14a_1(\ws_brp|dffe14a[1]~q ),
	.dffe14a_6(\ws_brp|dffe14a[6]~q ),
	.dffe14a_7(\ws_brp|dffe14a[7]~q ),
	.xor7(\ws_dgrp_gray2bin|xor7~combout ),
	.xor6(\ws_dgrp_gray2bin|xor6~combout ),
	.xor5(\ws_dgrp_gray2bin|xor5~combout ),
	.xor4(\ws_dgrp_gray2bin|xor4~combout ),
	.xor3(\ws_dgrp_gray2bin|xor3~combout ),
	.xor2(\ws_dgrp_gray2bin|xor2~combout ),
	.xor1(\ws_dgrp_gray2bin|xor1~combout ),
	.xor0(\ws_dgrp_gray2bin|xor0~combout ));

Computer_System_dffpipe_3dc_1 wraclr(
	.clock(wrclk),
	.dffe13a_0(dffe13a_0),
	.clrn(comb));

Computer_System_alt_synch_pipe_0ol rs_dgwp(
	.dffe17a_1(\rs_dgwp|dffpipe15|dffe17a[1]~q ),
	.dffe17a_6(\rs_dgwp|dffpipe15|dffe17a[6]~q ),
	.dffe17a_4(\rs_dgwp|dffpipe15|dffe17a[4]~q ),
	.dffe17a_5(\rs_dgwp|dffpipe15|dffe17a[5]~q ),
	.dffe17a_2(\rs_dgwp|dffpipe15|dffe17a[2]~q ),
	.dffe17a_3(\rs_dgwp|dffpipe15|dffe17a[3]~q ),
	.dffe17a_0(\rs_dgwp|dffpipe15|dffe17a[0]~q ),
	.dffe17a_8(\rs_dgwp|dffpipe15|dffe17a[8]~q ),
	.dffe17a_7(\rs_dgwp|dffpipe15|dffe17a[7]~q ),
	.clrn(\rdaclr|dffe13a[0]~q ),
	.delayed_wrptr_g_1(\delayed_wrptr_g[1]~q ),
	.delayed_wrptr_g_6(\delayed_wrptr_g[6]~q ),
	.delayed_wrptr_g_4(\delayed_wrptr_g[4]~q ),
	.delayed_wrptr_g_5(\delayed_wrptr_g[5]~q ),
	.delayed_wrptr_g_2(\delayed_wrptr_g[2]~q ),
	.delayed_wrptr_g_3(\delayed_wrptr_g[3]~q ),
	.delayed_wrptr_g_0(\delayed_wrptr_g[0]~q ),
	.delayed_wrptr_g_8(\delayed_wrptr_g[8]~q ),
	.delayed_wrptr_g_7(\delayed_wrptr_g[7]~q ),
	.clock(rdclk));

Computer_System_dffpipe_gd9_1 rs_bwp(
	.clrn(\rdaclr|dffe13a[0]~q ),
	.dffe14a_0(\rs_bwp|dffe14a[0]~q ),
	.dffe14a_1(\rs_bwp|dffe14a[1]~q ),
	.dffe14a_2(\rs_bwp|dffe14a[2]~q ),
	.dffe14a_3(\rs_bwp|dffe14a[3]~q ),
	.dffe14a_4(\rs_bwp|dffe14a[4]~q ),
	.dffe14a_5(\rs_bwp|dffe14a[5]~q ),
	.dffe14a_6(\rs_bwp|dffe14a[6]~q ),
	.dffe14a_7(\rs_bwp|dffe14a[7]~q ),
	.xor7(\rs_dgwp_gray2bin|xor7~combout ),
	.xor3(\rs_dgwp_gray2bin|xor3~combout ),
	.xor0(\rs_dgwp_gray2bin|xor0~combout ),
	.xor1(\rs_dgwp_gray2bin|xor1~combout ),
	.xor2(\rs_dgwp_gray2bin|xor2~combout ),
	.xor6(\rs_dgwp_gray2bin|xor6~combout ),
	.xor4(\rs_dgwp_gray2bin|xor4~combout ),
	.xor5(\rs_dgwp_gray2bin|xor5~combout ),
	.clock(rdclk));

Computer_System_dffpipe_gd9 rs_brp(
	.clrn(\rdaclr|dffe13a[0]~q ),
	.dffe14a_0(\rs_brp|dffe14a[0]~q ),
	.dffe14a_1(\rs_brp|dffe14a[1]~q ),
	.dffe14a_2(\rs_brp|dffe14a[2]~q ),
	.dffe14a_3(\rs_brp|dffe14a[3]~q ),
	.dffe14a_4(\rs_brp|dffe14a[4]~q ),
	.dffe14a_5(\rs_brp|dffe14a[5]~q ),
	.dffe14a_6(\rs_brp|dffe14a[6]~q ),
	.dffe14a_7(\rs_brp|dffe14a[7]~q ),
	.xor7(\rdptr_g_gray2bin|xor7~combout ),
	.xor3(\rdptr_g_gray2bin|xor3~combout ),
	.xor0(\rdptr_g_gray2bin|xor0~combout ),
	.xor1(\rdptr_g_gray2bin|xor1~combout ),
	.xor2(\rdptr_g_gray2bin|xor2~combout ),
	.xor6(\rdptr_g_gray2bin|xor6~combout ),
	.xor4(\rdptr_g_gray2bin|xor4~combout ),
	.xor5(\rdptr_g_gray2bin|xor5~combout ),
	.clock(rdclk));

Computer_System_dffpipe_3dc rdaclr(
	.dffe13a_0(\rdaclr|dffe13a[0]~q ),
	.clrn(comb),
	.clock(rdclk));

Computer_System_altsyncram_26d1 fifo_ram(
	.q_b({q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clock0(wrclk),
	.address_a({\ram_address_a[7]~combout ,\wrptr_g[6]~q ,\wrptr_g[5]~q ,\wrptr_g[4]~q ,\wrptr_g[3]~q ,\wrptr_g[2]~q ,wrptr_g_1,\wrptr_g[0]~q }),
	.wren_a(\wrptr_g1p|_~0_combout ),
	.aclr1(\rdaclr|dffe13a[0]~q ),
	.addressstall_b(\valid_rdreq~0_combout ),
	.clocken1(\valid_rdreq~0_combout ),
	.data_a({data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_b({\rdptr_g1p|_~0_combout ,\rdptr_g1p|counter5a6~q ,\rdptr_g1p|counter5a5~q ,\rdptr_g1p|counter5a4~q ,\rdptr_g1p|counter5a3~q ,\rdptr_g1p|counter5a2~q ,\rdptr_g1p|counter5a1~q ,\rdptr_g1p|counter5a0~_wirecell_combout }),
	.clock1(rdclk));

Computer_System_a_graycounter_bcc wrptr_g1p(
	.clock(wrclk),
	.op_2(op_23),
	.op_21(op_26),
	.op_22(op_27),
	.wrfull(wrfull),
	.wrfull1(wrfull1),
	.dffe13a_0(dffe13a_0),
	.wrfull2(wrfull2),
	.m0_write(m0_write),
	._(\wrptr_g1p|_~0_combout ),
	.wrfull3(wrfull3),
	.counter8a11(\wrptr_g1p|counter8a1~q ),
	.counter8a61(\wrptr_g1p|counter8a6~q ),
	.counter8a41(\wrptr_g1p|counter8a4~q ),
	.counter8a51(\wrptr_g1p|counter8a5~q ),
	.counter8a21(\wrptr_g1p|counter8a2~q ),
	.counter8a31(\wrptr_g1p|counter8a3~q ),
	.counter8a01(\wrptr_g1p|counter8a0~q ),
	.counter8a81(\wrptr_g1p|counter8a8~q ),
	.counter8a71(\wrptr_g1p|counter8a7~q ));

Computer_System_a_graycounter_fu6 rdptr_g1p(
	.aneb_result_wire_0(aneb_result_wire_03),
	.dffe13a_0(\rdaclr|dffe13a[0]~q ),
	.valid_rdreq(\valid_rdreq~0_combout ),
	.counter5a01(\rdptr_g1p|counter5a0~q ),
	.counter5a11(\rdptr_g1p|counter5a1~q ),
	.counter5a21(\rdptr_g1p|counter5a2~q ),
	.counter5a31(\rdptr_g1p|counter5a3~q ),
	.counter5a41(\rdptr_g1p|counter5a4~q ),
	.counter5a51(\rdptr_g1p|counter5a5~q ),
	.counter5a61(\rdptr_g1p|counter5a6~q ),
	.counter5a71(\rdptr_g1p|counter5a7~q ),
	.counter5a81(\rdptr_g1p|counter5a8~q ),
	._(\rdptr_g1p|_~0_combout ),
	.counter5a02(\rdptr_g1p|counter5a0~_wirecell_combout ),
	.fifo_hps_to_fpga_out_read(fifo_hps_to_fpga_out_read),
	.clock(rdclk));

Computer_System_a_gray2bin_g9b_3 ws_dgrp_gray2bin(
	.dffe20a_1(dffe20a_1),
	.dffe20a_6(\ws_dgrp|dffpipe18|dffe20a[6]~q ),
	.dffe20a_4(\ws_dgrp|dffpipe18|dffe20a[4]~q ),
	.dffe20a_5(\ws_dgrp|dffpipe18|dffe20a[5]~q ),
	.dffe20a_2(\ws_dgrp|dffpipe18|dffe20a[2]~q ),
	.dffe20a_3(\ws_dgrp|dffpipe18|dffe20a[3]~q ),
	.dffe20a_0(\ws_dgrp|dffpipe18|dffe20a[0]~q ),
	.dffe20a_8(\ws_dgrp|dffpipe18|dffe20a[8]~q ),
	.dffe20a_7(\ws_dgrp|dffpipe18|dffe20a[7]~q ),
	.xor71(\ws_dgrp_gray2bin|xor7~combout ),
	.xor61(\ws_dgrp_gray2bin|xor6~combout ),
	.xor51(\ws_dgrp_gray2bin|xor5~combout ),
	.xor41(\ws_dgrp_gray2bin|xor4~combout ),
	.xor31(\ws_dgrp_gray2bin|xor3~combout ),
	.xor21(\ws_dgrp_gray2bin|xor2~combout ),
	.xor11(\ws_dgrp_gray2bin|xor1~combout ),
	.xor01(\ws_dgrp_gray2bin|xor0~combout ));

Computer_System_a_gray2bin_g9b_2 wrptr_g_gray2bin(
	.wrptr_g_1(wrptr_g_1),
	.wrptr_g_6(\wrptr_g[6]~q ),
	.wrptr_g_4(\wrptr_g[4]~q ),
	.wrptr_g_5(\wrptr_g[5]~q ),
	.wrptr_g_2(\wrptr_g[2]~q ),
	.wrptr_g_3(\wrptr_g[3]~q ),
	.wrptr_g_0(\wrptr_g[0]~q ),
	.wrptr_g_8(\wrptr_g[8]~q ),
	.wrptr_g_7(\wrptr_g[7]~q ),
	.xor61(\wrptr_g_gray2bin|xor6~combout ),
	.xor51(\wrptr_g_gray2bin|xor5~combout ),
	.xor41(\wrptr_g_gray2bin|xor4~combout ),
	.xor31(\wrptr_g_gray2bin|xor3~combout ),
	.xor21(\wrptr_g_gray2bin|xor2~combout ),
	.xor11(\wrptr_g_gray2bin|xor1~combout ),
	.xor01(\wrptr_g_gray2bin|xor0~combout ));

Computer_System_a_gray2bin_g9b_1 rs_dgwp_gray2bin(
	.dffe17a_1(\rs_dgwp|dffpipe15|dffe17a[1]~q ),
	.dffe17a_6(\rs_dgwp|dffpipe15|dffe17a[6]~q ),
	.dffe17a_4(\rs_dgwp|dffpipe15|dffe17a[4]~q ),
	.dffe17a_5(\rs_dgwp|dffpipe15|dffe17a[5]~q ),
	.dffe17a_2(\rs_dgwp|dffpipe15|dffe17a[2]~q ),
	.dffe17a_3(\rs_dgwp|dffpipe15|dffe17a[3]~q ),
	.dffe17a_0(\rs_dgwp|dffpipe15|dffe17a[0]~q ),
	.dffe17a_8(\rs_dgwp|dffpipe15|dffe17a[8]~q ),
	.dffe17a_7(\rs_dgwp|dffpipe15|dffe17a[7]~q ),
	.xor71(\rs_dgwp_gray2bin|xor7~combout ),
	.xor31(\rs_dgwp_gray2bin|xor3~combout ),
	.xor01(\rs_dgwp_gray2bin|xor0~combout ),
	.xor11(\rs_dgwp_gray2bin|xor1~combout ),
	.xor21(\rs_dgwp_gray2bin|xor2~combout ),
	.xor61(\rs_dgwp_gray2bin|xor6~combout ),
	.xor41(\rs_dgwp_gray2bin|xor4~combout ),
	.xor51(\rs_dgwp_gray2bin|xor5~combout ));

Computer_System_a_gray2bin_g9b rdptr_g_gray2bin(
	.rdptr_g_1(\rdptr_g[1]~q ),
	.rdptr_g_6(\rdptr_g[6]~q ),
	.rdptr_g_4(\rdptr_g[4]~q ),
	.rdptr_g_5(\rdptr_g[5]~q ),
	.rdptr_g_2(\rdptr_g[2]~q ),
	.rdptr_g_3(\rdptr_g[3]~q ),
	.rdptr_g_0(\rdptr_g[0]~q ),
	.rdptr_g_8(\rdptr_g[8]~q ),
	.rdptr_g_7(\rdptr_g[7]~q ),
	.xor71(\rdptr_g_gray2bin|xor7~combout ),
	.xor31(\rdptr_g_gray2bin|xor3~combout ),
	.xor01(\rdptr_g_gray2bin|xor0~combout ),
	.xor11(\rdptr_g_gray2bin|xor1~combout ),
	.xor21(\rdptr_g_gray2bin|xor2~combout ),
	.xor61(\rdptr_g_gray2bin|xor6~combout ),
	.xor41(\rdptr_g_gray2bin|xor4~combout ),
	.xor51(\rdptr_g_gray2bin|xor5~combout ));

dffeas \rdptr_g[1] (
	.clk(rdclk),
	.d(\rdptr_g1p|counter5a1~q ),
	.asdata(vcc),
	.clrn(\rdaclr|dffe13a[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_rdreq~0_combout ),
	.q(\rdptr_g[1]~q ),
	.prn(vcc));
defparam \rdptr_g[1] .is_wysiwyg = "true";
defparam \rdptr_g[1] .power_up = "low";

dffeas \rdptr_g[6] (
	.clk(rdclk),
	.d(\rdptr_g1p|counter5a6~q ),
	.asdata(vcc),
	.clrn(\rdaclr|dffe13a[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_rdreq~0_combout ),
	.q(\rdptr_g[6]~q ),
	.prn(vcc));
defparam \rdptr_g[6] .is_wysiwyg = "true";
defparam \rdptr_g[6] .power_up = "low";

dffeas \rdptr_g[4] (
	.clk(rdclk),
	.d(\rdptr_g1p|counter5a4~q ),
	.asdata(vcc),
	.clrn(\rdaclr|dffe13a[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_rdreq~0_combout ),
	.q(\rdptr_g[4]~q ),
	.prn(vcc));
defparam \rdptr_g[4] .is_wysiwyg = "true";
defparam \rdptr_g[4] .power_up = "low";

dffeas \rdptr_g[5] (
	.clk(rdclk),
	.d(\rdptr_g1p|counter5a5~q ),
	.asdata(vcc),
	.clrn(\rdaclr|dffe13a[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_rdreq~0_combout ),
	.q(\rdptr_g[5]~q ),
	.prn(vcc));
defparam \rdptr_g[5] .is_wysiwyg = "true";
defparam \rdptr_g[5] .power_up = "low";

dffeas \rdptr_g[2] (
	.clk(rdclk),
	.d(\rdptr_g1p|counter5a2~q ),
	.asdata(vcc),
	.clrn(\rdaclr|dffe13a[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_rdreq~0_combout ),
	.q(\rdptr_g[2]~q ),
	.prn(vcc));
defparam \rdptr_g[2] .is_wysiwyg = "true";
defparam \rdptr_g[2] .power_up = "low";

dffeas \rdptr_g[3] (
	.clk(rdclk),
	.d(\rdptr_g1p|counter5a3~q ),
	.asdata(vcc),
	.clrn(\rdaclr|dffe13a[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_rdreq~0_combout ),
	.q(\rdptr_g[3]~q ),
	.prn(vcc));
defparam \rdptr_g[3] .is_wysiwyg = "true";
defparam \rdptr_g[3] .power_up = "low";

dffeas \rdptr_g[0] (
	.clk(rdclk),
	.d(\rdptr_g[0]~0_combout ),
	.asdata(vcc),
	.clrn(\rdaclr|dffe13a[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_rdreq~0_combout ),
	.q(\rdptr_g[0]~q ),
	.prn(vcc));
defparam \rdptr_g[0] .is_wysiwyg = "true";
defparam \rdptr_g[0] .power_up = "low";

dffeas \rdptr_g[8] (
	.clk(rdclk),
	.d(\rdptr_g1p|counter5a8~q ),
	.asdata(vcc),
	.clrn(\rdaclr|dffe13a[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_rdreq~0_combout ),
	.q(\rdptr_g[8]~q ),
	.prn(vcc));
defparam \rdptr_g[8] .is_wysiwyg = "true";
defparam \rdptr_g[8] .power_up = "low";

dffeas \rdptr_g[7] (
	.clk(rdclk),
	.d(\rdptr_g1p|counter5a7~q ),
	.asdata(vcc),
	.clrn(\rdaclr|dffe13a[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_rdreq~0_combout ),
	.q(\rdptr_g[7]~q ),
	.prn(vcc));
defparam \rdptr_g[7] .is_wysiwyg = "true";
defparam \rdptr_g[7] .power_up = "low";

dffeas \wrptr_g[6] (
	.clk(wrclk),
	.d(\wrptr_g1p|counter8a6~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wrptr_g1p|_~0_combout ),
	.q(\wrptr_g[6]~q ),
	.prn(vcc));
defparam \wrptr_g[6] .is_wysiwyg = "true";
defparam \wrptr_g[6] .power_up = "low";

dffeas \wrptr_g[4] (
	.clk(wrclk),
	.d(\wrptr_g1p|counter8a4~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wrptr_g1p|_~0_combout ),
	.q(\wrptr_g[4]~q ),
	.prn(vcc));
defparam \wrptr_g[4] .is_wysiwyg = "true";
defparam \wrptr_g[4] .power_up = "low";

dffeas \wrptr_g[5] (
	.clk(wrclk),
	.d(\wrptr_g1p|counter8a5~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wrptr_g1p|_~0_combout ),
	.q(\wrptr_g[5]~q ),
	.prn(vcc));
defparam \wrptr_g[5] .is_wysiwyg = "true";
defparam \wrptr_g[5] .power_up = "low";

dffeas \wrptr_g[2] (
	.clk(wrclk),
	.d(\wrptr_g1p|counter8a2~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wrptr_g1p|_~0_combout ),
	.q(\wrptr_g[2]~q ),
	.prn(vcc));
defparam \wrptr_g[2] .is_wysiwyg = "true";
defparam \wrptr_g[2] .power_up = "low";

dffeas \wrptr_g[3] (
	.clk(wrclk),
	.d(\wrptr_g1p|counter8a3~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wrptr_g1p|_~0_combout ),
	.q(\wrptr_g[3]~q ),
	.prn(vcc));
defparam \wrptr_g[3] .is_wysiwyg = "true";
defparam \wrptr_g[3] .power_up = "low";

dffeas \wrptr_g[0] (
	.clk(wrclk),
	.d(\wrptr_g[0]~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wrptr_g1p|_~0_combout ),
	.q(\wrptr_g[0]~q ),
	.prn(vcc));
defparam \wrptr_g[0] .is_wysiwyg = "true";
defparam \wrptr_g[0] .power_up = "low";

dffeas \wrptr_g[8] (
	.clk(wrclk),
	.d(\wrptr_g1p|counter8a8~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wrptr_g1p|_~0_combout ),
	.q(\wrptr_g[8]~q ),
	.prn(vcc));
defparam \wrptr_g[8] .is_wysiwyg = "true";
defparam \wrptr_g[8] .power_up = "low";

dffeas \wrptr_g[7] (
	.clk(wrclk),
	.d(\wrptr_g1p|counter8a7~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wrptr_g1p|_~0_combout ),
	.q(\wrptr_g[7]~q ),
	.prn(vcc));
defparam \wrptr_g[7] .is_wysiwyg = "true";
defparam \wrptr_g[7] .power_up = "low";

cyclonev_lcell_comb \valid_rdreq~0 (
	.dataa(!data_wire_2),
	.datab(!fifo_hps_to_fpga_out_read),
	.datac(!\rdaclr|dffe13a[0]~q ),
	.datad(!aneb_result_wire_0),
	.datae(!aneb_result_wire_01),
	.dataf(!aneb_result_wire_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\valid_rdreq~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \valid_rdreq~0 .extended_lut = "off";
defparam \valid_rdreq~0 .lut_mask = 64'h0303030303030301;
defparam \valid_rdreq~0 .shared_arith = "off";

cyclonev_lcell_comb \ram_address_a[7] (
	.dataa(!\wrptr_g[8]~q ),
	.datab(!\wrptr_g[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_address_a[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_address_a[7] .extended_lut = "off";
defparam \ram_address_a[7] .lut_mask = 64'h6666666666666666;
defparam \ram_address_a[7] .shared_arith = "off";

dffeas \delayed_wrptr_g[1] (
	.clk(wrclk),
	.d(wrptr_g_1),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_wrptr_g[1]~q ),
	.prn(vcc));
defparam \delayed_wrptr_g[1] .is_wysiwyg = "true";
defparam \delayed_wrptr_g[1] .power_up = "low";

dffeas \delayed_wrptr_g[6] (
	.clk(wrclk),
	.d(\wrptr_g[6]~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_wrptr_g[6]~q ),
	.prn(vcc));
defparam \delayed_wrptr_g[6] .is_wysiwyg = "true";
defparam \delayed_wrptr_g[6] .power_up = "low";

dffeas \delayed_wrptr_g[4] (
	.clk(wrclk),
	.d(\wrptr_g[4]~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_wrptr_g[4]~q ),
	.prn(vcc));
defparam \delayed_wrptr_g[4] .is_wysiwyg = "true";
defparam \delayed_wrptr_g[4] .power_up = "low";

dffeas \delayed_wrptr_g[5] (
	.clk(wrclk),
	.d(\wrptr_g[5]~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_wrptr_g[5]~q ),
	.prn(vcc));
defparam \delayed_wrptr_g[5] .is_wysiwyg = "true";
defparam \delayed_wrptr_g[5] .power_up = "low";

dffeas \delayed_wrptr_g[2] (
	.clk(wrclk),
	.d(\wrptr_g[2]~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_wrptr_g[2]~q ),
	.prn(vcc));
defparam \delayed_wrptr_g[2] .is_wysiwyg = "true";
defparam \delayed_wrptr_g[2] .power_up = "low";

dffeas \delayed_wrptr_g[3] (
	.clk(wrclk),
	.d(\wrptr_g[3]~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_wrptr_g[3]~q ),
	.prn(vcc));
defparam \delayed_wrptr_g[3] .is_wysiwyg = "true";
defparam \delayed_wrptr_g[3] .power_up = "low";

dffeas \delayed_wrptr_g[0] (
	.clk(wrclk),
	.d(\wrptr_g[0]~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_wrptr_g[0]~q ),
	.prn(vcc));
defparam \delayed_wrptr_g[0] .is_wysiwyg = "true";
defparam \delayed_wrptr_g[0] .power_up = "low";

dffeas \delayed_wrptr_g[8] (
	.clk(wrclk),
	.d(\wrptr_g[8]~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_wrptr_g[8]~q ),
	.prn(vcc));
defparam \delayed_wrptr_g[8] .is_wysiwyg = "true";
defparam \delayed_wrptr_g[8] .power_up = "low";

dffeas \delayed_wrptr_g[7] (
	.clk(wrclk),
	.d(\wrptr_g[7]~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_wrptr_g[7]~q ),
	.prn(vcc));
defparam \delayed_wrptr_g[7] .is_wysiwyg = "true";
defparam \delayed_wrptr_g[7] .power_up = "low";

cyclonev_lcell_comb \rdptr_g[0]~0 (
	.dataa(!\rdptr_g1p|counter5a0~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdptr_g[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdptr_g[0]~0 .extended_lut = "off";
defparam \rdptr_g[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdptr_g[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \wrptr_g[0]~0 (
	.dataa(!\wrptr_g1p|counter8a0~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wrptr_g[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wrptr_g[0]~0 .extended_lut = "off";
defparam \wrptr_g[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wrptr_g[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \op_2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\ws_brp|dffe14a[2]~q ),
	.datad(!\ws_bwp|dffe14a[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_2~22 ),
	.sharein(\op_2~23 ),
	.combout(),
	.sumout(op_2),
	.cout(\op_2~2 ),
	.shareout(\op_2~3 ));
defparam \op_2~1 .extended_lut = "off";
defparam \op_2~1 .lut_mask = 64'h000000F00000F00F;
defparam \op_2~1 .shared_arith = "on";

cyclonev_lcell_comb \op_2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\ws_brp|dffe14a[3]~q ),
	.datad(!\ws_bwp|dffe14a[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_2~2 ),
	.sharein(\op_2~3 ),
	.combout(),
	.sumout(op_21),
	.cout(\op_2~6 ),
	.shareout(\op_2~7 ));
defparam \op_2~5 .extended_lut = "off";
defparam \op_2~5 .lut_mask = 64'h000000F00000F00F;
defparam \op_2~5 .shared_arith = "on";

cyclonev_lcell_comb \op_2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\ws_brp|dffe14a[4]~q ),
	.datad(!\ws_bwp|dffe14a[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_2~6 ),
	.sharein(\op_2~7 ),
	.combout(),
	.sumout(op_22),
	.cout(\op_2~10 ),
	.shareout(\op_2~11 ));
defparam \op_2~9 .extended_lut = "off";
defparam \op_2~9 .lut_mask = 64'h000000F00000F00F;
defparam \op_2~9 .shared_arith = "on";

cyclonev_lcell_comb \op_2~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\ws_brp|dffe14a[5]~q ),
	.datad(!\ws_bwp|dffe14a[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_2~10 ),
	.sharein(\op_2~11 ),
	.combout(),
	.sumout(op_23),
	.cout(\op_2~14 ),
	.shareout(\op_2~15 ));
defparam \op_2~13 .extended_lut = "off";
defparam \op_2~13 .lut_mask = 64'h000000F00000F00F;
defparam \op_2~13 .shared_arith = "on";

cyclonev_lcell_comb \op_2~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\ws_brp|dffe14a[0]~q ),
	.datad(!\ws_bwp|dffe14a[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(op_24),
	.cout(\op_2~18 ),
	.shareout(\op_2~19 ));
defparam \op_2~17 .extended_lut = "off";
defparam \op_2~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \op_2~17 .shared_arith = "on";

cyclonev_lcell_comb \op_2~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\ws_brp|dffe14a[1]~q ),
	.datad(!\ws_bwp|dffe14a[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_2~18 ),
	.sharein(\op_2~19 ),
	.combout(),
	.sumout(op_25),
	.cout(\op_2~22 ),
	.shareout(\op_2~23 ));
defparam \op_2~21 .extended_lut = "off";
defparam \op_2~21 .lut_mask = 64'h000000F00000F00F;
defparam \op_2~21 .shared_arith = "on";

cyclonev_lcell_comb \op_2~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\ws_brp|dffe14a[6]~q ),
	.datad(!\ws_bwp|dffe14a[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_2~14 ),
	.sharein(\op_2~15 ),
	.combout(),
	.sumout(op_26),
	.cout(\op_2~26 ),
	.shareout(\op_2~27 ));
defparam \op_2~25 .extended_lut = "off";
defparam \op_2~25 .lut_mask = 64'h000000F00000F00F;
defparam \op_2~25 .shared_arith = "on";

cyclonev_lcell_comb \op_2~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\ws_brp|dffe14a[7]~q ),
	.datad(!\ws_bwp|dffe14a[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_2~26 ),
	.sharein(\op_2~27 ),
	.combout(),
	.sumout(op_27),
	.cout(),
	.shareout());
defparam \op_2~29 .extended_lut = "off";
defparam \op_2~29 .lut_mask = 64'h000000000000F00F;
defparam \op_2~29 .shared_arith = "on";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rs_brp|dffe14a[0]~q ),
	.datad(!\rs_bwp|dffe14a[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(op_1),
	.cout(\op_1~2 ),
	.shareout(\op_1~3 ));
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \op_1~1 .shared_arith = "on";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rs_brp|dffe14a[1]~q ),
	.datad(!\rs_bwp|dffe14a[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(\op_1~3 ),
	.combout(),
	.sumout(op_11),
	.cout(\op_1~6 ),
	.shareout(\op_1~7 ));
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h000000F00000F00F;
defparam \op_1~5 .shared_arith = "on";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rs_brp|dffe14a[2]~q ),
	.datad(!\rs_bwp|dffe14a[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(\op_1~7 ),
	.combout(),
	.sumout(op_12),
	.cout(\op_1~10 ),
	.shareout(\op_1~11 ));
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h000000F00000F00F;
defparam \op_1~9 .shared_arith = "on";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rs_brp|dffe14a[3]~q ),
	.datad(!\rs_bwp|dffe14a[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(\op_1~11 ),
	.combout(),
	.sumout(op_13),
	.cout(\op_1~14 ),
	.shareout(\op_1~15 ));
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h000000F00000F00F;
defparam \op_1~13 .shared_arith = "on";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rs_brp|dffe14a[4]~q ),
	.datad(!\rs_bwp|dffe14a[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(\op_1~15 ),
	.combout(),
	.sumout(op_14),
	.cout(\op_1~18 ),
	.shareout(\op_1~19 ));
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h000000F00000F00F;
defparam \op_1~17 .shared_arith = "on";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rs_brp|dffe14a[5]~q ),
	.datad(!\rs_bwp|dffe14a[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(\op_1~19 ),
	.combout(),
	.sumout(op_15),
	.cout(\op_1~22 ),
	.shareout(\op_1~23 ));
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h000000F00000F00F;
defparam \op_1~21 .shared_arith = "on";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rs_brp|dffe14a[6]~q ),
	.datad(!\rs_bwp|dffe14a[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(\op_1~23 ),
	.combout(),
	.sumout(op_16),
	.cout(\op_1~26 ),
	.shareout(\op_1~27 ));
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h000000F00000F00F;
defparam \op_1~25 .shared_arith = "on";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rs_brp|dffe14a[7]~q ),
	.datad(!\rs_bwp|dffe14a[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(\op_1~27 ),
	.combout(),
	.sumout(op_17),
	.cout(),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h000000000000F00F;
defparam \op_1~29 .shared_arith = "on";

dffeas \wrptr_g[1] (
	.clk(wrclk),
	.d(\wrptr_g1p|counter8a1~q ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wrptr_g1p|_~0_combout ),
	.q(wrptr_g_1),
	.prn(vcc));
defparam \wrptr_g[1] .is_wysiwyg = "true";
defparam \wrptr_g[1] .power_up = "low";

endmodule

module Computer_System_a_gray2bin_g9b (
	rdptr_g_1,
	rdptr_g_6,
	rdptr_g_4,
	rdptr_g_5,
	rdptr_g_2,
	rdptr_g_3,
	rdptr_g_0,
	rdptr_g_8,
	rdptr_g_7,
	xor71,
	xor31,
	xor01,
	xor11,
	xor21,
	xor61,
	xor41,
	xor51)/* synthesis synthesis_greybox=0 */;
input 	rdptr_g_1;
input 	rdptr_g_6;
input 	rdptr_g_4;
input 	rdptr_g_5;
input 	rdptr_g_2;
input 	rdptr_g_3;
input 	rdptr_g_0;
input 	rdptr_g_8;
input 	rdptr_g_7;
output 	xor71;
output 	xor31;
output 	xor01;
output 	xor11;
output 	xor21;
output 	xor61;
output 	xor41;
output 	xor51;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb xor7(
	.dataa(!rdptr_g_8),
	.datab(!rdptr_g_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor71),
	.sumout(),
	.cout(),
	.shareout());
defparam xor7.extended_lut = "off";
defparam xor7.lut_mask = 64'h6666666666666666;
defparam xor7.shared_arith = "off";

cyclonev_lcell_comb xor3(
	.dataa(!rdptr_g_6),
	.datab(!rdptr_g_4),
	.datac(!rdptr_g_5),
	.datad(!rdptr_g_3),
	.datae(!xor71),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor31),
	.sumout(),
	.cout(),
	.shareout());
defparam xor3.extended_lut = "off";
defparam xor3.lut_mask = 64'h6996966969969669;
defparam xor3.shared_arith = "off";

cyclonev_lcell_comb xor0(
	.dataa(!rdptr_g_2),
	.datab(!rdptr_g_0),
	.datac(!rdptr_g_1),
	.datad(!xor31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor01),
	.sumout(),
	.cout(),
	.shareout());
defparam xor0.extended_lut = "off";
defparam xor0.lut_mask = 64'h6996699669966996;
defparam xor0.shared_arith = "off";

cyclonev_lcell_comb xor1(
	.dataa(!rdptr_g_2),
	.datab(!rdptr_g_1),
	.datac(!xor31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor11),
	.sumout(),
	.cout(),
	.shareout());
defparam xor1.extended_lut = "off";
defparam xor1.lut_mask = 64'h6969696969696969;
defparam xor1.shared_arith = "off";

cyclonev_lcell_comb xor2(
	.dataa(!rdptr_g_2),
	.datab(!xor31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor21),
	.sumout(),
	.cout(),
	.shareout());
defparam xor2.extended_lut = "off";
defparam xor2.lut_mask = 64'h6666666666666666;
defparam xor2.shared_arith = "off";

cyclonev_lcell_comb xor6(
	.dataa(!rdptr_g_6),
	.datab(!xor71),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor61),
	.sumout(),
	.cout(),
	.shareout());
defparam xor6.extended_lut = "off";
defparam xor6.lut_mask = 64'h6666666666666666;
defparam xor6.shared_arith = "off";

cyclonev_lcell_comb xor4(
	.dataa(!rdptr_g_4),
	.datab(!rdptr_g_5),
	.datac(!xor61),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor41),
	.sumout(),
	.cout(),
	.shareout());
defparam xor4.extended_lut = "off";
defparam xor4.lut_mask = 64'h6969696969696969;
defparam xor4.shared_arith = "off";

cyclonev_lcell_comb xor5(
	.dataa(!rdptr_g_5),
	.datab(!xor61),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor51),
	.sumout(),
	.cout(),
	.shareout());
defparam xor5.extended_lut = "off";
defparam xor5.lut_mask = 64'h6666666666666666;
defparam xor5.shared_arith = "off";

endmodule

module Computer_System_a_gray2bin_g9b_1 (
	dffe17a_1,
	dffe17a_6,
	dffe17a_4,
	dffe17a_5,
	dffe17a_2,
	dffe17a_3,
	dffe17a_0,
	dffe17a_8,
	dffe17a_7,
	xor71,
	xor31,
	xor01,
	xor11,
	xor21,
	xor61,
	xor41,
	xor51)/* synthesis synthesis_greybox=0 */;
input 	dffe17a_1;
input 	dffe17a_6;
input 	dffe17a_4;
input 	dffe17a_5;
input 	dffe17a_2;
input 	dffe17a_3;
input 	dffe17a_0;
input 	dffe17a_8;
input 	dffe17a_7;
output 	xor71;
output 	xor31;
output 	xor01;
output 	xor11;
output 	xor21;
output 	xor61;
output 	xor41;
output 	xor51;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb xor7(
	.dataa(!dffe17a_8),
	.datab(!dffe17a_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor71),
	.sumout(),
	.cout(),
	.shareout());
defparam xor7.extended_lut = "off";
defparam xor7.lut_mask = 64'h6666666666666666;
defparam xor7.shared_arith = "off";

cyclonev_lcell_comb xor3(
	.dataa(!dffe17a_6),
	.datab(!dffe17a_4),
	.datac(!dffe17a_5),
	.datad(!dffe17a_3),
	.datae(!xor71),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor31),
	.sumout(),
	.cout(),
	.shareout());
defparam xor3.extended_lut = "off";
defparam xor3.lut_mask = 64'h6996966969969669;
defparam xor3.shared_arith = "off";

cyclonev_lcell_comb xor0(
	.dataa(!dffe17a_2),
	.datab(!dffe17a_0),
	.datac(!dffe17a_1),
	.datad(!xor31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor01),
	.sumout(),
	.cout(),
	.shareout());
defparam xor0.extended_lut = "off";
defparam xor0.lut_mask = 64'h6996699669966996;
defparam xor0.shared_arith = "off";

cyclonev_lcell_comb xor1(
	.dataa(!dffe17a_2),
	.datab(!dffe17a_1),
	.datac(!xor31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor11),
	.sumout(),
	.cout(),
	.shareout());
defparam xor1.extended_lut = "off";
defparam xor1.lut_mask = 64'h6969696969696969;
defparam xor1.shared_arith = "off";

cyclonev_lcell_comb xor2(
	.dataa(!dffe17a_2),
	.datab(!xor31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor21),
	.sumout(),
	.cout(),
	.shareout());
defparam xor2.extended_lut = "off";
defparam xor2.lut_mask = 64'h6666666666666666;
defparam xor2.shared_arith = "off";

cyclonev_lcell_comb xor6(
	.dataa(!dffe17a_6),
	.datab(!xor71),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor61),
	.sumout(),
	.cout(),
	.shareout());
defparam xor6.extended_lut = "off";
defparam xor6.lut_mask = 64'h6666666666666666;
defparam xor6.shared_arith = "off";

cyclonev_lcell_comb xor4(
	.dataa(!dffe17a_4),
	.datab(!dffe17a_5),
	.datac(!xor61),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor41),
	.sumout(),
	.cout(),
	.shareout());
defparam xor4.extended_lut = "off";
defparam xor4.lut_mask = 64'h6969696969696969;
defparam xor4.shared_arith = "off";

cyclonev_lcell_comb xor5(
	.dataa(!dffe17a_5),
	.datab(!xor61),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor51),
	.sumout(),
	.cout(),
	.shareout());
defparam xor5.extended_lut = "off";
defparam xor5.lut_mask = 64'h6666666666666666;
defparam xor5.shared_arith = "off";

endmodule

module Computer_System_a_gray2bin_g9b_2 (
	wrptr_g_1,
	wrptr_g_6,
	wrptr_g_4,
	wrptr_g_5,
	wrptr_g_2,
	wrptr_g_3,
	wrptr_g_0,
	wrptr_g_8,
	wrptr_g_7,
	xor61,
	xor51,
	xor41,
	xor31,
	xor21,
	xor11,
	xor01)/* synthesis synthesis_greybox=0 */;
input 	wrptr_g_1;
input 	wrptr_g_6;
input 	wrptr_g_4;
input 	wrptr_g_5;
input 	wrptr_g_2;
input 	wrptr_g_3;
input 	wrptr_g_0;
input 	wrptr_g_8;
input 	wrptr_g_7;
output 	xor61;
output 	xor51;
output 	xor41;
output 	xor31;
output 	xor21;
output 	xor11;
output 	xor01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb xor6(
	.dataa(!wrptr_g_6),
	.datab(!wrptr_g_8),
	.datac(!wrptr_g_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor61),
	.sumout(),
	.cout(),
	.shareout());
defparam xor6.extended_lut = "off";
defparam xor6.lut_mask = 64'h6969696969696969;
defparam xor6.shared_arith = "off";

cyclonev_lcell_comb xor5(
	.dataa(!wrptr_g_5),
	.datab(!xor61),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor51),
	.sumout(),
	.cout(),
	.shareout());
defparam xor5.extended_lut = "off";
defparam xor5.lut_mask = 64'h6666666666666666;
defparam xor5.shared_arith = "off";

cyclonev_lcell_comb xor4(
	.dataa(!wrptr_g_4),
	.datab(!wrptr_g_5),
	.datac(!xor61),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor41),
	.sumout(),
	.cout(),
	.shareout());
defparam xor4.extended_lut = "off";
defparam xor4.lut_mask = 64'h6969696969696969;
defparam xor4.shared_arith = "off";

cyclonev_lcell_comb xor3(
	.dataa(!wrptr_g_3),
	.datab(!xor41),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor31),
	.sumout(),
	.cout(),
	.shareout());
defparam xor3.extended_lut = "off";
defparam xor3.lut_mask = 64'h6666666666666666;
defparam xor3.shared_arith = "off";

cyclonev_lcell_comb xor2(
	.dataa(!wrptr_g_2),
	.datab(!xor31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor21),
	.sumout(),
	.cout(),
	.shareout());
defparam xor2.extended_lut = "off";
defparam xor2.lut_mask = 64'h6666666666666666;
defparam xor2.shared_arith = "off";

cyclonev_lcell_comb xor1(
	.dataa(!wrptr_g_1),
	.datab(!xor21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor11),
	.sumout(),
	.cout(),
	.shareout());
defparam xor1.extended_lut = "off";
defparam xor1.lut_mask = 64'h6666666666666666;
defparam xor1.shared_arith = "off";

cyclonev_lcell_comb xor0(
	.dataa(!wrptr_g_0),
	.datab(!xor11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor01),
	.sumout(),
	.cout(),
	.shareout());
defparam xor0.extended_lut = "off";
defparam xor0.lut_mask = 64'h6666666666666666;
defparam xor0.shared_arith = "off";

endmodule

module Computer_System_a_gray2bin_g9b_3 (
	dffe20a_1,
	dffe20a_6,
	dffe20a_4,
	dffe20a_5,
	dffe20a_2,
	dffe20a_3,
	dffe20a_0,
	dffe20a_8,
	dffe20a_7,
	xor71,
	xor61,
	xor51,
	xor41,
	xor31,
	xor21,
	xor11,
	xor01)/* synthesis synthesis_greybox=0 */;
input 	dffe20a_1;
input 	dffe20a_6;
input 	dffe20a_4;
input 	dffe20a_5;
input 	dffe20a_2;
input 	dffe20a_3;
input 	dffe20a_0;
input 	dffe20a_8;
input 	dffe20a_7;
output 	xor71;
output 	xor61;
output 	xor51;
output 	xor41;
output 	xor31;
output 	xor21;
output 	xor11;
output 	xor01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb xor7(
	.dataa(!dffe20a_8),
	.datab(!dffe20a_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor71),
	.sumout(),
	.cout(),
	.shareout());
defparam xor7.extended_lut = "off";
defparam xor7.lut_mask = 64'h6666666666666666;
defparam xor7.shared_arith = "off";

cyclonev_lcell_comb xor6(
	.dataa(!dffe20a_6),
	.datab(!dffe20a_8),
	.datac(!dffe20a_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor61),
	.sumout(),
	.cout(),
	.shareout());
defparam xor6.extended_lut = "off";
defparam xor6.lut_mask = 64'h6969696969696969;
defparam xor6.shared_arith = "off";

cyclonev_lcell_comb xor5(
	.dataa(!dffe20a_5),
	.datab(!xor61),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor51),
	.sumout(),
	.cout(),
	.shareout());
defparam xor5.extended_lut = "off";
defparam xor5.lut_mask = 64'h6666666666666666;
defparam xor5.shared_arith = "off";

cyclonev_lcell_comb xor4(
	.dataa(!dffe20a_4),
	.datab(!dffe20a_5),
	.datac(!xor61),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor41),
	.sumout(),
	.cout(),
	.shareout());
defparam xor4.extended_lut = "off";
defparam xor4.lut_mask = 64'h6969696969696969;
defparam xor4.shared_arith = "off";

cyclonev_lcell_comb xor3(
	.dataa(!dffe20a_3),
	.datab(!xor41),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor31),
	.sumout(),
	.cout(),
	.shareout());
defparam xor3.extended_lut = "off";
defparam xor3.lut_mask = 64'h6666666666666666;
defparam xor3.shared_arith = "off";

cyclonev_lcell_comb xor2(
	.dataa(!dffe20a_2),
	.datab(!xor31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor21),
	.sumout(),
	.cout(),
	.shareout());
defparam xor2.extended_lut = "off";
defparam xor2.lut_mask = 64'h6666666666666666;
defparam xor2.shared_arith = "off";

cyclonev_lcell_comb xor1(
	.dataa(!dffe20a_1),
	.datab(!xor21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor11),
	.sumout(),
	.cout(),
	.shareout());
defparam xor1.extended_lut = "off";
defparam xor1.lut_mask = 64'h6666666666666666;
defparam xor1.shared_arith = "off";

cyclonev_lcell_comb xor0(
	.dataa(!dffe20a_0),
	.datab(!xor11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xor01),
	.sumout(),
	.cout(),
	.shareout());
defparam xor0.extended_lut = "off";
defparam xor0.lut_mask = 64'h6666666666666666;
defparam xor0.shared_arith = "off";

endmodule

module Computer_System_a_graycounter_bcc (
	clock,
	op_2,
	op_21,
	op_22,
	wrfull,
	wrfull1,
	dffe13a_0,
	wrfull2,
	m0_write,
	_,
	wrfull3,
	counter8a11,
	counter8a61,
	counter8a41,
	counter8a51,
	counter8a21,
	counter8a31,
	counter8a01,
	counter8a81,
	counter8a71)/* synthesis synthesis_greybox=0 */;
input 	clock;
input 	op_2;
input 	op_21;
input 	op_22;
input 	wrfull;
input 	wrfull1;
input 	dffe13a_0;
input 	wrfull2;
input 	m0_write;
output 	_;
input 	wrfull3;
output 	counter8a11;
output 	counter8a61;
output 	counter8a41;
output 	counter8a51;
output 	counter8a21;
output 	counter8a31;
output 	counter8a01;
output 	counter8a81;
output 	counter8a71;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~3_combout ;
wire \sub_parity10a[1]~q ;
wire \_~4_combout ;
wire \sub_parity10a[0]~q ;
wire \_~2_combout ;
wire \parity9~q ;
wire \counter8a1~0_combout ;
wire \cntr_cout[2]~1_combout ;
wire \cntr_cout[2]~0_combout ;
wire \counter8a6~0_combout ;
wire \counter8a4~0_combout ;
wire \counter8a5~0_combout ;
wire \counter8a2~0_combout ;
wire \counter8a3~0_combout ;
wire \counter8a0~0_combout ;
wire \_~1_combout ;
wire \counter8a8~0_combout ;
wire \counter8a7~0_combout ;


cyclonev_lcell_comb \_~0 (
	.dataa(!wrfull2),
	.datab(!m0_write),
	.datac(!op_21),
	.datad(!op_22),
	.datae(!op_2),
	.dataf(!wrfull3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(_),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'h1111111111111110;
defparam \_~0 .shared_arith = "off";

dffeas counter8a1(
	.clk(clock),
	.d(\counter8a1~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter8a11),
	.prn(vcc));
defparam counter8a1.is_wysiwyg = "true";
defparam counter8a1.power_up = "low";

dffeas counter8a6(
	.clk(clock),
	.d(\counter8a6~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter8a61),
	.prn(vcc));
defparam counter8a6.is_wysiwyg = "true";
defparam counter8a6.power_up = "low";

dffeas counter8a4(
	.clk(clock),
	.d(\counter8a4~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter8a41),
	.prn(vcc));
defparam counter8a4.is_wysiwyg = "true";
defparam counter8a4.power_up = "low";

dffeas counter8a5(
	.clk(clock),
	.d(\counter8a5~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter8a51),
	.prn(vcc));
defparam counter8a5.is_wysiwyg = "true";
defparam counter8a5.power_up = "low";

dffeas counter8a2(
	.clk(clock),
	.d(\counter8a2~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter8a21),
	.prn(vcc));
defparam counter8a2.is_wysiwyg = "true";
defparam counter8a2.power_up = "low";

dffeas counter8a3(
	.clk(clock),
	.d(\counter8a3~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter8a31),
	.prn(vcc));
defparam counter8a3.is_wysiwyg = "true";
defparam counter8a3.power_up = "low";

dffeas counter8a0(
	.clk(clock),
	.d(\counter8a0~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter8a01),
	.prn(vcc));
defparam counter8a0.is_wysiwyg = "true";
defparam counter8a0.power_up = "low";

dffeas counter8a8(
	.clk(clock),
	.d(\counter8a8~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter8a81),
	.prn(vcc));
defparam counter8a8.is_wysiwyg = "true";
defparam counter8a8.power_up = "low";

dffeas counter8a7(
	.clk(clock),
	.d(\counter8a7~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter8a71),
	.prn(vcc));
defparam counter8a7.is_wysiwyg = "true";
defparam counter8a7.power_up = "low";

cyclonev_lcell_comb \_~3 (
	.dataa(!counter8a81),
	.datab(!counter8a71),
	.datac(!counter8a61),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~3 .extended_lut = "off";
defparam \_~3 .lut_mask = 64'h6969696969696969;
defparam \_~3 .shared_arith = "off";

dffeas \sub_parity10a[1] (
	.clk(clock),
	.d(\_~3_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(\sub_parity10a[1]~q ),
	.prn(vcc));
defparam \sub_parity10a[1] .is_wysiwyg = "true";
defparam \sub_parity10a[1] .power_up = "low";

cyclonev_lcell_comb \_~4 (
	.dataa(!counter8a41),
	.datab(!counter8a51),
	.datac(!counter8a21),
	.datad(!counter8a31),
	.datae(!counter8a01),
	.dataf(!counter8a11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~4 .extended_lut = "off";
defparam \_~4 .lut_mask = 64'h9669699669969669;
defparam \_~4 .shared_arith = "off";

dffeas \sub_parity10a[0] (
	.clk(clock),
	.d(\_~4_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(\sub_parity10a[0]~q ),
	.prn(vcc));
defparam \sub_parity10a[0] .is_wysiwyg = "true";
defparam \sub_parity10a[0] .power_up = "low";

cyclonev_lcell_comb \_~2 (
	.dataa(!\sub_parity10a[1]~q ),
	.datab(!\sub_parity10a[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~2 .extended_lut = "off";
defparam \_~2 .lut_mask = 64'h9999999999999999;
defparam \_~2 .shared_arith = "off";

dffeas parity9(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(\parity9~q ),
	.prn(vcc));
defparam parity9.is_wysiwyg = "true";
defparam parity9.power_up = "low";

cyclonev_lcell_comb \counter8a1~0 (
	.dataa(!_),
	.datab(!counter8a01),
	.datac(!counter8a11),
	.datad(!\parity9~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter8a1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter8a1~0 .extended_lut = "off";
defparam \counter8a1~0 .lut_mask = 64'h4B0F4B0F4B0F4B0F;
defparam \counter8a1~0 .shared_arith = "off";

cyclonev_lcell_comb \cntr_cout[2]~1 (
	.dataa(!counter8a11),
	.datab(!\parity9~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cntr_cout[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cntr_cout[2]~1 .extended_lut = "off";
defparam \cntr_cout[2]~1 .lut_mask = 64'h8888888888888888;
defparam \cntr_cout[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \cntr_cout[2]~0 (
	.dataa(!counter8a01),
	.datab(!wrfull),
	.datac(!wrfull1),
	.datad(!wrfull2),
	.datae(!m0_write),
	.dataf(!\cntr_cout[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cntr_cout[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cntr_cout[2]~0 .extended_lut = "off";
defparam \cntr_cout[2]~0 .lut_mask = 64'h0000000000000054;
defparam \cntr_cout[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \counter8a6~0 (
	.dataa(!counter8a61),
	.datab(!counter8a51),
	.datac(!counter8a41),
	.datad(!counter8a21),
	.datae(!counter8a31),
	.dataf(!\cntr_cout[2]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter8a6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter8a6~0 .extended_lut = "off";
defparam \counter8a6~0 .lut_mask = 64'h5555555565555555;
defparam \counter8a6~0 .shared_arith = "off";

cyclonev_lcell_comb \counter8a4~0 (
	.dataa(!counter8a41),
	.datab(!counter8a21),
	.datac(!counter8a31),
	.datad(!\cntr_cout[2]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter8a4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter8a4~0 .extended_lut = "off";
defparam \counter8a4~0 .lut_mask = 64'h5559555955595559;
defparam \counter8a4~0 .shared_arith = "off";

cyclonev_lcell_comb \counter8a5~0 (
	.dataa(!counter8a41),
	.datab(!counter8a51),
	.datac(!counter8a21),
	.datad(!counter8a31),
	.datae(!\cntr_cout[2]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter8a5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter8a5~0 .extended_lut = "off";
defparam \counter8a5~0 .lut_mask = 64'h3333633333336333;
defparam \counter8a5~0 .shared_arith = "off";

cyclonev_lcell_comb \counter8a2~0 (
	.dataa(!_),
	.datab(!counter8a21),
	.datac(!counter8a01),
	.datad(!counter8a11),
	.datae(!\parity9~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter8a2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter8a2~0 .extended_lut = "off";
defparam \counter8a2~0 .lut_mask = 64'h3336333333363333;
defparam \counter8a2~0 .shared_arith = "off";

cyclonev_lcell_comb \counter8a3~0 (
	.dataa(!counter8a21),
	.datab(!counter8a31),
	.datac(!\cntr_cout[2]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter8a3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter8a3~0 .extended_lut = "off";
defparam \counter8a3~0 .lut_mask = 64'h3636363636363636;
defparam \counter8a3~0 .shared_arith = "off";

cyclonev_lcell_comb \counter8a0~0 (
	.dataa(!_),
	.datab(!counter8a01),
	.datac(!\parity9~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter8a0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter8a0~0 .extended_lut = "off";
defparam \counter8a0~0 .lut_mask = 64'h3636363636363636;
defparam \counter8a0~0 .shared_arith = "off";

cyclonev_lcell_comb \_~1 (
	.dataa(!counter8a41),
	.datab(!counter8a21),
	.datac(!counter8a31),
	.datad(!\cntr_cout[2]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~1 .extended_lut = "off";
defparam \_~1 .lut_mask = 64'h0080008000800080;
defparam \_~1 .shared_arith = "off";

cyclonev_lcell_comb \counter8a8~0 (
	.dataa(!counter8a81),
	.datab(!counter8a61),
	.datac(!counter8a51),
	.datad(!\_~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter8a8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter8a8~0 .extended_lut = "off";
defparam \counter8a8~0 .lut_mask = 64'h5595559555955595;
defparam \counter8a8~0 .shared_arith = "off";

cyclonev_lcell_comb \counter8a7~0 (
	.dataa(!counter8a71),
	.datab(!counter8a61),
	.datac(!counter8a51),
	.datad(!\_~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter8a7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter8a7~0 .extended_lut = "off";
defparam \counter8a7~0 .lut_mask = 64'h5565556555655565;
defparam \counter8a7~0 .shared_arith = "off";

endmodule

module Computer_System_a_graycounter_fu6 (
	aneb_result_wire_0,
	dffe13a_0,
	valid_rdreq,
	counter5a01,
	counter5a11,
	counter5a21,
	counter5a31,
	counter5a41,
	counter5a51,
	counter5a61,
	counter5a71,
	counter5a81,
	_,
	counter5a02,
	fifo_hps_to_fpga_out_read,
	clock)/* synthesis synthesis_greybox=0 */;
input 	aneb_result_wire_0;
input 	dffe13a_0;
input 	valid_rdreq;
output 	counter5a01;
output 	counter5a11;
output 	counter5a21;
output 	counter5a31;
output 	counter5a41;
output 	counter5a51;
output 	counter5a61;
output 	counter5a71;
output 	counter5a81;
output 	_;
output 	counter5a02;
input 	fifo_hps_to_fpga_out_read;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~4_combout ;
wire \sub_parity7a[1]~q ;
wire \_~5_combout ;
wire \sub_parity7a[0]~q ;
wire \_~3_combout ;
wire \parity6~q ;
wire \counter5a0~0_combout ;
wire \counter5a1~0_combout ;
wire \counter5a2~0_combout ;
wire \counter5a3~0_combout ;
wire \_~1_combout ;
wire \counter5a4~0_combout ;
wire \counter5a5~0_combout ;
wire \counter5a6~0_combout ;
wire \_~2_combout ;
wire \counter5a7~0_combout ;
wire \counter5a8~0_combout ;


dffeas counter5a0(
	.clk(clock),
	.d(\counter5a0~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter5a01),
	.prn(vcc));
defparam counter5a0.is_wysiwyg = "true";
defparam counter5a0.power_up = "low";

dffeas counter5a1(
	.clk(clock),
	.d(\counter5a1~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter5a11),
	.prn(vcc));
defparam counter5a1.is_wysiwyg = "true";
defparam counter5a1.power_up = "low";

dffeas counter5a2(
	.clk(clock),
	.d(\counter5a2~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter5a21),
	.prn(vcc));
defparam counter5a2.is_wysiwyg = "true";
defparam counter5a2.power_up = "low";

dffeas counter5a3(
	.clk(clock),
	.d(\counter5a3~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter5a31),
	.prn(vcc));
defparam counter5a3.is_wysiwyg = "true";
defparam counter5a3.power_up = "low";

dffeas counter5a4(
	.clk(clock),
	.d(\counter5a4~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter5a41),
	.prn(vcc));
defparam counter5a4.is_wysiwyg = "true";
defparam counter5a4.power_up = "low";

dffeas counter5a5(
	.clk(clock),
	.d(\counter5a5~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter5a51),
	.prn(vcc));
defparam counter5a5.is_wysiwyg = "true";
defparam counter5a5.power_up = "low";

dffeas counter5a6(
	.clk(clock),
	.d(\counter5a6~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter5a61),
	.prn(vcc));
defparam counter5a6.is_wysiwyg = "true";
defparam counter5a6.power_up = "low";

dffeas counter5a7(
	.clk(clock),
	.d(\counter5a7~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter5a71),
	.prn(vcc));
defparam counter5a7.is_wysiwyg = "true";
defparam counter5a7.power_up = "low";

dffeas counter5a8(
	.clk(clock),
	.d(\counter5a8~0_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(counter5a81),
	.prn(vcc));
defparam counter5a8.is_wysiwyg = "true";
defparam counter5a8.power_up = "low";

cyclonev_lcell_comb \_~0 (
	.dataa(!counter5a71),
	.datab(!counter5a81),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(_),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'h6666666666666666;
defparam \_~0 .shared_arith = "off";

cyclonev_lcell_comb \counter5a0~_wirecell (
	.dataa(!counter5a01),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(counter5a02),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter5a0~_wirecell .extended_lut = "off";
defparam \counter5a0~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter5a0~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \_~4 (
	.dataa(!counter5a61),
	.datab(!_),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~4 .extended_lut = "off";
defparam \_~4 .lut_mask = 64'h6666666666666666;
defparam \_~4 .shared_arith = "off";

dffeas \sub_parity7a[1] (
	.clk(clock),
	.d(\_~4_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(valid_rdreq),
	.q(\sub_parity7a[1]~q ),
	.prn(vcc));
defparam \sub_parity7a[1] .is_wysiwyg = "true";
defparam \sub_parity7a[1] .power_up = "low";

cyclonev_lcell_comb \_~5 (
	.dataa(!counter5a01),
	.datab(!counter5a11),
	.datac(!counter5a21),
	.datad(!counter5a31),
	.datae(!counter5a41),
	.dataf(!counter5a51),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~5 .extended_lut = "off";
defparam \_~5 .lut_mask = 64'h9669699669969669;
defparam \_~5 .shared_arith = "off";

dffeas \sub_parity7a[0] (
	.clk(clock),
	.d(\_~5_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(valid_rdreq),
	.q(\sub_parity7a[0]~q ),
	.prn(vcc));
defparam \sub_parity7a[0] .is_wysiwyg = "true";
defparam \sub_parity7a[0] .power_up = "low";

cyclonev_lcell_comb \_~3 (
	.dataa(!\sub_parity7a[1]~q ),
	.datab(!\sub_parity7a[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~3 .extended_lut = "off";
defparam \_~3 .lut_mask = 64'h9999999999999999;
defparam \_~3 .shared_arith = "off";

dffeas parity6(
	.clk(clock),
	.d(\_~3_combout ),
	.asdata(vcc),
	.clrn(dffe13a_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(valid_rdreq),
	.q(\parity6~q ),
	.prn(vcc));
defparam parity6.is_wysiwyg = "true";
defparam parity6.power_up = "low";

cyclonev_lcell_comb \counter5a0~0 (
	.dataa(!fifo_hps_to_fpga_out_read),
	.datab(!dffe13a_0),
	.datac(!counter5a01),
	.datad(!\parity6~q ),
	.datae(!aneb_result_wire_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter5a0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter5a0~0 .extended_lut = "off";
defparam \counter5a0~0 .lut_mask = 64'h0F0F0F1E0F0F0F1E;
defparam \counter5a0~0 .shared_arith = "off";

cyclonev_lcell_comb \counter5a1~0 (
	.dataa(!fifo_hps_to_fpga_out_read),
	.datab(!dffe13a_0),
	.datac(!counter5a01),
	.datad(!counter5a11),
	.datae(!\parity6~q ),
	.dataf(!aneb_result_wire_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter5a1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter5a1~0 .extended_lut = "off";
defparam \counter5a1~0 .lut_mask = 64'h00FF00FF10EF00FF;
defparam \counter5a1~0 .shared_arith = "off";

cyclonev_lcell_comb \counter5a2~0 (
	.dataa(!counter5a01),
	.datab(!counter5a11),
	.datac(!counter5a21),
	.datad(!\parity6~q ),
	.datae(!valid_rdreq),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter5a2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter5a2~0 .extended_lut = "off";
defparam \counter5a2~0 .lut_mask = 64'h0F0F1E0F0F0F1E0F;
defparam \counter5a2~0 .shared_arith = "off";

cyclonev_lcell_comb \counter5a3~0 (
	.dataa(!counter5a01),
	.datab(!counter5a11),
	.datac(!counter5a21),
	.datad(!counter5a31),
	.datae(!\parity6~q ),
	.dataf(!valid_rdreq),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter5a3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter5a3~0 .extended_lut = "off";
defparam \counter5a3~0 .lut_mask = 64'h00FF00FF04FB00FF;
defparam \counter5a3~0 .shared_arith = "off";

cyclonev_lcell_comb \_~1 (
	.dataa(!fifo_hps_to_fpga_out_read),
	.datab(!dffe13a_0),
	.datac(!counter5a01),
	.datad(!counter5a11),
	.datae(!\parity6~q ),
	.dataf(!aneb_result_wire_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~1 .extended_lut = "off";
defparam \_~1 .lut_mask = 64'h0000000001000000;
defparam \_~1 .shared_arith = "off";

cyclonev_lcell_comb \counter5a4~0 (
	.dataa(!counter5a21),
	.datab(!counter5a31),
	.datac(!counter5a41),
	.datad(!\_~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter5a4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter5a4~0 .extended_lut = "off";
defparam \counter5a4~0 .lut_mask = 64'h0F2D0F2D0F2D0F2D;
defparam \counter5a4~0 .shared_arith = "off";

cyclonev_lcell_comb \counter5a5~0 (
	.dataa(!counter5a21),
	.datab(!counter5a31),
	.datac(!counter5a41),
	.datad(!counter5a51),
	.datae(!\_~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter5a5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter5a5~0 .extended_lut = "off";
defparam \counter5a5~0 .lut_mask = 64'h00FF08F700FF08F7;
defparam \counter5a5~0 .shared_arith = "off";

cyclonev_lcell_comb \counter5a6~0 (
	.dataa(!counter5a21),
	.datab(!counter5a31),
	.datac(!counter5a41),
	.datad(!counter5a51),
	.datae(!counter5a61),
	.dataf(!\_~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter5a6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter5a6~0 .extended_lut = "off";
defparam \counter5a6~0 .lut_mask = 64'h0000FFFF0080FF7F;
defparam \counter5a6~0 .shared_arith = "off";

cyclonev_lcell_comb \_~2 (
	.dataa(!counter5a01),
	.datab(!counter5a11),
	.datac(!counter5a21),
	.datad(!\parity6~q ),
	.datae(!valid_rdreq),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~2 .extended_lut = "off";
defparam \_~2 .lut_mask = 64'h0000400000004000;
defparam \_~2 .shared_arith = "off";

cyclonev_lcell_comb \counter5a7~0 (
	.dataa(!counter5a31),
	.datab(!counter5a41),
	.datac(!counter5a51),
	.datad(!counter5a61),
	.datae(!counter5a71),
	.dataf(!\_~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter5a7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter5a7~0 .extended_lut = "off";
defparam \counter5a7~0 .lut_mask = 64'h0000FFFF0080FF7F;
defparam \counter5a7~0 .shared_arith = "off";

cyclonev_lcell_comb \counter5a8~0 (
	.dataa(!counter5a31),
	.datab(!counter5a41),
	.datac(!counter5a51),
	.datad(!counter5a61),
	.datae(!counter5a81),
	.dataf(!\_~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter5a8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter5a8~0 .extended_lut = "off";
defparam \counter5a8~0 .lut_mask = 64'h0000FFFF80007FFF;
defparam \counter5a8~0 .shared_arith = "off";

endmodule

module Computer_System_alt_synch_pipe_0ol (
	dffe17a_1,
	dffe17a_6,
	dffe17a_4,
	dffe17a_5,
	dffe17a_2,
	dffe17a_3,
	dffe17a_0,
	dffe17a_8,
	dffe17a_7,
	clrn,
	delayed_wrptr_g_1,
	delayed_wrptr_g_6,
	delayed_wrptr_g_4,
	delayed_wrptr_g_5,
	delayed_wrptr_g_2,
	delayed_wrptr_g_3,
	delayed_wrptr_g_0,
	delayed_wrptr_g_8,
	delayed_wrptr_g_7,
	clock)/* synthesis synthesis_greybox=0 */;
output 	dffe17a_1;
output 	dffe17a_6;
output 	dffe17a_4;
output 	dffe17a_5;
output 	dffe17a_2;
output 	dffe17a_3;
output 	dffe17a_0;
output 	dffe17a_8;
output 	dffe17a_7;
input 	clrn;
input 	delayed_wrptr_g_1;
input 	delayed_wrptr_g_6;
input 	delayed_wrptr_g_4;
input 	delayed_wrptr_g_5;
input 	delayed_wrptr_g_2;
input 	delayed_wrptr_g_3;
input 	delayed_wrptr_g_0;
input 	delayed_wrptr_g_8;
input 	delayed_wrptr_g_7;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_dffpipe_hd9 dffpipe15(
	.dffe17a_1(dffe17a_1),
	.dffe17a_6(dffe17a_6),
	.dffe17a_4(dffe17a_4),
	.dffe17a_5(dffe17a_5),
	.dffe17a_2(dffe17a_2),
	.dffe17a_3(dffe17a_3),
	.dffe17a_0(dffe17a_0),
	.dffe17a_8(dffe17a_8),
	.dffe17a_7(dffe17a_7),
	.clrn(clrn),
	.delayed_wrptr_g_1(delayed_wrptr_g_1),
	.delayed_wrptr_g_6(delayed_wrptr_g_6),
	.delayed_wrptr_g_4(delayed_wrptr_g_4),
	.delayed_wrptr_g_5(delayed_wrptr_g_5),
	.delayed_wrptr_g_2(delayed_wrptr_g_2),
	.delayed_wrptr_g_3(delayed_wrptr_g_3),
	.delayed_wrptr_g_0(delayed_wrptr_g_0),
	.delayed_wrptr_g_8(delayed_wrptr_g_8),
	.delayed_wrptr_g_7(delayed_wrptr_g_7),
	.clock(clock));

endmodule

module Computer_System_dffpipe_hd9 (
	dffe17a_1,
	dffe17a_6,
	dffe17a_4,
	dffe17a_5,
	dffe17a_2,
	dffe17a_3,
	dffe17a_0,
	dffe17a_8,
	dffe17a_7,
	clrn,
	delayed_wrptr_g_1,
	delayed_wrptr_g_6,
	delayed_wrptr_g_4,
	delayed_wrptr_g_5,
	delayed_wrptr_g_2,
	delayed_wrptr_g_3,
	delayed_wrptr_g_0,
	delayed_wrptr_g_8,
	delayed_wrptr_g_7,
	clock)/* synthesis synthesis_greybox=0 */;
output 	dffe17a_1;
output 	dffe17a_6;
output 	dffe17a_4;
output 	dffe17a_5;
output 	dffe17a_2;
output 	dffe17a_3;
output 	dffe17a_0;
output 	dffe17a_8;
output 	dffe17a_7;
input 	clrn;
input 	delayed_wrptr_g_1;
input 	delayed_wrptr_g_6;
input 	delayed_wrptr_g_4;
input 	delayed_wrptr_g_5;
input 	delayed_wrptr_g_2;
input 	delayed_wrptr_g_3;
input 	delayed_wrptr_g_0;
input 	delayed_wrptr_g_8;
input 	delayed_wrptr_g_7;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffe16a[1]~q ;
wire \dffe16a[6]~q ;
wire \dffe16a[4]~q ;
wire \dffe16a[5]~q ;
wire \dffe16a[2]~q ;
wire \dffe16a[3]~q ;
wire \dffe16a[0]~q ;
wire \dffe16a[8]~q ;
wire \dffe16a[7]~q ;


dffeas \dffe17a[1] (
	.clk(clock),
	.d(\dffe16a[1]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe17a_1),
	.prn(vcc));
defparam \dffe17a[1] .is_wysiwyg = "true";
defparam \dffe17a[1] .power_up = "low";
defparam \dffe17a[1] .x_on_violation = "off";

dffeas \dffe17a[6] (
	.clk(clock),
	.d(\dffe16a[6]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe17a_6),
	.prn(vcc));
defparam \dffe17a[6] .is_wysiwyg = "true";
defparam \dffe17a[6] .power_up = "low";
defparam \dffe17a[6] .x_on_violation = "off";

dffeas \dffe17a[4] (
	.clk(clock),
	.d(\dffe16a[4]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe17a_4),
	.prn(vcc));
defparam \dffe17a[4] .is_wysiwyg = "true";
defparam \dffe17a[4] .power_up = "low";
defparam \dffe17a[4] .x_on_violation = "off";

dffeas \dffe17a[5] (
	.clk(clock),
	.d(\dffe16a[5]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe17a_5),
	.prn(vcc));
defparam \dffe17a[5] .is_wysiwyg = "true";
defparam \dffe17a[5] .power_up = "low";
defparam \dffe17a[5] .x_on_violation = "off";

dffeas \dffe17a[2] (
	.clk(clock),
	.d(\dffe16a[2]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe17a_2),
	.prn(vcc));
defparam \dffe17a[2] .is_wysiwyg = "true";
defparam \dffe17a[2] .power_up = "low";
defparam \dffe17a[2] .x_on_violation = "off";

dffeas \dffe17a[3] (
	.clk(clock),
	.d(\dffe16a[3]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe17a_3),
	.prn(vcc));
defparam \dffe17a[3] .is_wysiwyg = "true";
defparam \dffe17a[3] .power_up = "low";
defparam \dffe17a[3] .x_on_violation = "off";

dffeas \dffe17a[0] (
	.clk(clock),
	.d(\dffe16a[0]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe17a_0),
	.prn(vcc));
defparam \dffe17a[0] .is_wysiwyg = "true";
defparam \dffe17a[0] .power_up = "low";
defparam \dffe17a[0] .x_on_violation = "off";

dffeas \dffe17a[8] (
	.clk(clock),
	.d(\dffe16a[8]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe17a_8),
	.prn(vcc));
defparam \dffe17a[8] .is_wysiwyg = "true";
defparam \dffe17a[8] .power_up = "low";
defparam \dffe17a[8] .x_on_violation = "off";

dffeas \dffe17a[7] (
	.clk(clock),
	.d(\dffe16a[7]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe17a_7),
	.prn(vcc));
defparam \dffe17a[7] .is_wysiwyg = "true";
defparam \dffe17a[7] .power_up = "low";
defparam \dffe17a[7] .x_on_violation = "off";

dffeas \dffe16a[1] (
	.clk(clock),
	.d(delayed_wrptr_g_1),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe16a[1]~q ),
	.prn(vcc));
defparam \dffe16a[1] .is_wysiwyg = "true";
defparam \dffe16a[1] .power_up = "low";
defparam \dffe16a[1] .x_on_violation = "off";

dffeas \dffe16a[6] (
	.clk(clock),
	.d(delayed_wrptr_g_6),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe16a[6]~q ),
	.prn(vcc));
defparam \dffe16a[6] .is_wysiwyg = "true";
defparam \dffe16a[6] .power_up = "low";
defparam \dffe16a[6] .x_on_violation = "off";

dffeas \dffe16a[4] (
	.clk(clock),
	.d(delayed_wrptr_g_4),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe16a[4]~q ),
	.prn(vcc));
defparam \dffe16a[4] .is_wysiwyg = "true";
defparam \dffe16a[4] .power_up = "low";
defparam \dffe16a[4] .x_on_violation = "off";

dffeas \dffe16a[5] (
	.clk(clock),
	.d(delayed_wrptr_g_5),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe16a[5]~q ),
	.prn(vcc));
defparam \dffe16a[5] .is_wysiwyg = "true";
defparam \dffe16a[5] .power_up = "low";
defparam \dffe16a[5] .x_on_violation = "off";

dffeas \dffe16a[2] (
	.clk(clock),
	.d(delayed_wrptr_g_2),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe16a[2]~q ),
	.prn(vcc));
defparam \dffe16a[2] .is_wysiwyg = "true";
defparam \dffe16a[2] .power_up = "low";
defparam \dffe16a[2] .x_on_violation = "off";

dffeas \dffe16a[3] (
	.clk(clock),
	.d(delayed_wrptr_g_3),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe16a[3]~q ),
	.prn(vcc));
defparam \dffe16a[3] .is_wysiwyg = "true";
defparam \dffe16a[3] .power_up = "low";
defparam \dffe16a[3] .x_on_violation = "off";

dffeas \dffe16a[0] (
	.clk(clock),
	.d(delayed_wrptr_g_0),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe16a[0]~q ),
	.prn(vcc));
defparam \dffe16a[0] .is_wysiwyg = "true";
defparam \dffe16a[0] .power_up = "low";
defparam \dffe16a[0] .x_on_violation = "off";

dffeas \dffe16a[8] (
	.clk(clock),
	.d(delayed_wrptr_g_8),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe16a[8]~q ),
	.prn(vcc));
defparam \dffe16a[8] .is_wysiwyg = "true";
defparam \dffe16a[8] .power_up = "low";
defparam \dffe16a[8] .x_on_violation = "off";

dffeas \dffe16a[7] (
	.clk(clock),
	.d(delayed_wrptr_g_7),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe16a[7]~q ),
	.prn(vcc));
defparam \dffe16a[7] .is_wysiwyg = "true";
defparam \dffe16a[7] .power_up = "low";
defparam \dffe16a[7] .x_on_violation = "off";

endmodule

module Computer_System_alt_synch_pipe_1ol (
	clock,
	rdptr_g_1,
	rdptr_g_6,
	rdptr_g_4,
	rdptr_g_5,
	rdptr_g_2,
	rdptr_g_3,
	rdptr_g_0,
	rdptr_g_8,
	rdptr_g_7,
	clrn,
	dffe20a_1,
	dffe20a_6,
	dffe20a_4,
	dffe20a_5,
	dffe20a_2,
	dffe20a_3,
	dffe20a_0,
	dffe20a_8,
	dffe20a_7)/* synthesis synthesis_greybox=0 */;
input 	clock;
input 	rdptr_g_1;
input 	rdptr_g_6;
input 	rdptr_g_4;
input 	rdptr_g_5;
input 	rdptr_g_2;
input 	rdptr_g_3;
input 	rdptr_g_0;
input 	rdptr_g_8;
input 	rdptr_g_7;
input 	clrn;
output 	dffe20a_1;
output 	dffe20a_6;
output 	dffe20a_4;
output 	dffe20a_5;
output 	dffe20a_2;
output 	dffe20a_3;
output 	dffe20a_0;
output 	dffe20a_8;
output 	dffe20a_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_dffpipe_id9 dffpipe18(
	.clock(clock),
	.rdptr_g_1(rdptr_g_1),
	.rdptr_g_6(rdptr_g_6),
	.rdptr_g_4(rdptr_g_4),
	.rdptr_g_5(rdptr_g_5),
	.rdptr_g_2(rdptr_g_2),
	.rdptr_g_3(rdptr_g_3),
	.rdptr_g_0(rdptr_g_0),
	.rdptr_g_8(rdptr_g_8),
	.rdptr_g_7(rdptr_g_7),
	.clrn(clrn),
	.dffe20a_1(dffe20a_1),
	.dffe20a_6(dffe20a_6),
	.dffe20a_4(dffe20a_4),
	.dffe20a_5(dffe20a_5),
	.dffe20a_2(dffe20a_2),
	.dffe20a_3(dffe20a_3),
	.dffe20a_0(dffe20a_0),
	.dffe20a_8(dffe20a_8),
	.dffe20a_7(dffe20a_7));

endmodule

module Computer_System_dffpipe_id9 (
	clock,
	rdptr_g_1,
	rdptr_g_6,
	rdptr_g_4,
	rdptr_g_5,
	rdptr_g_2,
	rdptr_g_3,
	rdptr_g_0,
	rdptr_g_8,
	rdptr_g_7,
	clrn,
	dffe20a_1,
	dffe20a_6,
	dffe20a_4,
	dffe20a_5,
	dffe20a_2,
	dffe20a_3,
	dffe20a_0,
	dffe20a_8,
	dffe20a_7)/* synthesis synthesis_greybox=0 */;
input 	clock;
input 	rdptr_g_1;
input 	rdptr_g_6;
input 	rdptr_g_4;
input 	rdptr_g_5;
input 	rdptr_g_2;
input 	rdptr_g_3;
input 	rdptr_g_0;
input 	rdptr_g_8;
input 	rdptr_g_7;
input 	clrn;
output 	dffe20a_1;
output 	dffe20a_6;
output 	dffe20a_4;
output 	dffe20a_5;
output 	dffe20a_2;
output 	dffe20a_3;
output 	dffe20a_0;
output 	dffe20a_8;
output 	dffe20a_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffe19a[1]~q ;
wire \dffe19a[6]~q ;
wire \dffe19a[4]~q ;
wire \dffe19a[5]~q ;
wire \dffe19a[2]~q ;
wire \dffe19a[3]~q ;
wire \dffe19a[0]~q ;
wire \dffe19a[8]~q ;
wire \dffe19a[7]~q ;


dffeas \dffe20a[1] (
	.clk(clock),
	.d(\dffe19a[1]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe20a_1),
	.prn(vcc));
defparam \dffe20a[1] .is_wysiwyg = "true";
defparam \dffe20a[1] .power_up = "low";
defparam \dffe20a[1] .x_on_violation = "off";

dffeas \dffe20a[6] (
	.clk(clock),
	.d(\dffe19a[6]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe20a_6),
	.prn(vcc));
defparam \dffe20a[6] .is_wysiwyg = "true";
defparam \dffe20a[6] .power_up = "low";
defparam \dffe20a[6] .x_on_violation = "off";

dffeas \dffe20a[4] (
	.clk(clock),
	.d(\dffe19a[4]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe20a_4),
	.prn(vcc));
defparam \dffe20a[4] .is_wysiwyg = "true";
defparam \dffe20a[4] .power_up = "low";
defparam \dffe20a[4] .x_on_violation = "off";

dffeas \dffe20a[5] (
	.clk(clock),
	.d(\dffe19a[5]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe20a_5),
	.prn(vcc));
defparam \dffe20a[5] .is_wysiwyg = "true";
defparam \dffe20a[5] .power_up = "low";
defparam \dffe20a[5] .x_on_violation = "off";

dffeas \dffe20a[2] (
	.clk(clock),
	.d(\dffe19a[2]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe20a_2),
	.prn(vcc));
defparam \dffe20a[2] .is_wysiwyg = "true";
defparam \dffe20a[2] .power_up = "low";
defparam \dffe20a[2] .x_on_violation = "off";

dffeas \dffe20a[3] (
	.clk(clock),
	.d(\dffe19a[3]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe20a_3),
	.prn(vcc));
defparam \dffe20a[3] .is_wysiwyg = "true";
defparam \dffe20a[3] .power_up = "low";
defparam \dffe20a[3] .x_on_violation = "off";

dffeas \dffe20a[0] (
	.clk(clock),
	.d(\dffe19a[0]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe20a_0),
	.prn(vcc));
defparam \dffe20a[0] .is_wysiwyg = "true";
defparam \dffe20a[0] .power_up = "low";
defparam \dffe20a[0] .x_on_violation = "off";

dffeas \dffe20a[8] (
	.clk(clock),
	.d(\dffe19a[8]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe20a_8),
	.prn(vcc));
defparam \dffe20a[8] .is_wysiwyg = "true";
defparam \dffe20a[8] .power_up = "low";
defparam \dffe20a[8] .x_on_violation = "off";

dffeas \dffe20a[7] (
	.clk(clock),
	.d(\dffe19a[7]~q ),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe20a_7),
	.prn(vcc));
defparam \dffe20a[7] .is_wysiwyg = "true";
defparam \dffe20a[7] .power_up = "low";
defparam \dffe20a[7] .x_on_violation = "off";

dffeas \dffe19a[1] (
	.clk(clock),
	.d(rdptr_g_1),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe19a[1]~q ),
	.prn(vcc));
defparam \dffe19a[1] .is_wysiwyg = "true";
defparam \dffe19a[1] .power_up = "low";
defparam \dffe19a[1] .x_on_violation = "off";

dffeas \dffe19a[6] (
	.clk(clock),
	.d(rdptr_g_6),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe19a[6]~q ),
	.prn(vcc));
defparam \dffe19a[6] .is_wysiwyg = "true";
defparam \dffe19a[6] .power_up = "low";
defparam \dffe19a[6] .x_on_violation = "off";

dffeas \dffe19a[4] (
	.clk(clock),
	.d(rdptr_g_4),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe19a[4]~q ),
	.prn(vcc));
defparam \dffe19a[4] .is_wysiwyg = "true";
defparam \dffe19a[4] .power_up = "low";
defparam \dffe19a[4] .x_on_violation = "off";

dffeas \dffe19a[5] (
	.clk(clock),
	.d(rdptr_g_5),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe19a[5]~q ),
	.prn(vcc));
defparam \dffe19a[5] .is_wysiwyg = "true";
defparam \dffe19a[5] .power_up = "low";
defparam \dffe19a[5] .x_on_violation = "off";

dffeas \dffe19a[2] (
	.clk(clock),
	.d(rdptr_g_2),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe19a[2]~q ),
	.prn(vcc));
defparam \dffe19a[2] .is_wysiwyg = "true";
defparam \dffe19a[2] .power_up = "low";
defparam \dffe19a[2] .x_on_violation = "off";

dffeas \dffe19a[3] (
	.clk(clock),
	.d(rdptr_g_3),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe19a[3]~q ),
	.prn(vcc));
defparam \dffe19a[3] .is_wysiwyg = "true";
defparam \dffe19a[3] .power_up = "low";
defparam \dffe19a[3] .x_on_violation = "off";

dffeas \dffe19a[0] (
	.clk(clock),
	.d(rdptr_g_0),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe19a[0]~q ),
	.prn(vcc));
defparam \dffe19a[0] .is_wysiwyg = "true";
defparam \dffe19a[0] .power_up = "low";
defparam \dffe19a[0] .x_on_violation = "off";

dffeas \dffe19a[8] (
	.clk(clock),
	.d(rdptr_g_8),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe19a[8]~q ),
	.prn(vcc));
defparam \dffe19a[8] .is_wysiwyg = "true";
defparam \dffe19a[8] .power_up = "low";
defparam \dffe19a[8] .x_on_violation = "off";

dffeas \dffe19a[7] (
	.clk(clock),
	.d(rdptr_g_7),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe19a[7]~q ),
	.prn(vcc));
defparam \dffe19a[7] .is_wysiwyg = "true";
defparam \dffe19a[7] .power_up = "low";
defparam \dffe19a[7] .x_on_violation = "off";

endmodule

module Computer_System_altsyncram_26d1 (
	q_b,
	clock0,
	address_a,
	wren_a,
	aclr1,
	addressstall_b,
	clocken1,
	data_a,
	address_b,
	clock1)/* synthesis synthesis_greybox=0 */;
output 	[31:0] q_b;
input 	clock0;
input 	[7:0] address_a;
input 	wren_a;
input 	aclr1;
input 	addressstall_b;
input 	clocken1;
input 	[31:0] data_a;
input 	[7:0] address_b;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block11a0_PORTBDATAOUT_bus;
wire [143:0] ram_block11a1_PORTBDATAOUT_bus;
wire [143:0] ram_block11a2_PORTBDATAOUT_bus;
wire [143:0] ram_block11a3_PORTBDATAOUT_bus;
wire [143:0] ram_block11a4_PORTBDATAOUT_bus;
wire [143:0] ram_block11a5_PORTBDATAOUT_bus;
wire [143:0] ram_block11a6_PORTBDATAOUT_bus;
wire [143:0] ram_block11a7_PORTBDATAOUT_bus;
wire [143:0] ram_block11a8_PORTBDATAOUT_bus;
wire [143:0] ram_block11a9_PORTBDATAOUT_bus;
wire [143:0] ram_block11a10_PORTBDATAOUT_bus;
wire [143:0] ram_block11a11_PORTBDATAOUT_bus;
wire [143:0] ram_block11a12_PORTBDATAOUT_bus;
wire [143:0] ram_block11a13_PORTBDATAOUT_bus;
wire [143:0] ram_block11a14_PORTBDATAOUT_bus;
wire [143:0] ram_block11a15_PORTBDATAOUT_bus;
wire [143:0] ram_block11a16_PORTBDATAOUT_bus;
wire [143:0] ram_block11a17_PORTBDATAOUT_bus;
wire [143:0] ram_block11a18_PORTBDATAOUT_bus;
wire [143:0] ram_block11a19_PORTBDATAOUT_bus;
wire [143:0] ram_block11a20_PORTBDATAOUT_bus;
wire [143:0] ram_block11a21_PORTBDATAOUT_bus;
wire [143:0] ram_block11a22_PORTBDATAOUT_bus;
wire [143:0] ram_block11a23_PORTBDATAOUT_bus;
wire [143:0] ram_block11a24_PORTBDATAOUT_bus;
wire [143:0] ram_block11a25_PORTBDATAOUT_bus;
wire [143:0] ram_block11a26_PORTBDATAOUT_bus;
wire [143:0] ram_block11a27_PORTBDATAOUT_bus;
wire [143:0] ram_block11a28_PORTBDATAOUT_bus;
wire [143:0] ram_block11a29_PORTBDATAOUT_bus;
wire [143:0] ram_block11a30_PORTBDATAOUT_bus;
wire [143:0] ram_block11a31_PORTBDATAOUT_bus;

assign q_b[0] = ram_block11a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block11a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block11a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block11a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block11a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block11a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block11a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block11a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block11a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block11a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block11a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block11a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block11a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block11a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block11a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block11a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block11a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block11a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block11a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block11a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block11a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block11a21_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block11a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block11a23_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block11a24_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block11a25_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block11a26_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block11a27_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block11a28_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block11a29_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block11a30_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block11a31_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block11a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a0.clk0_core_clock_enable = "ena0";
defparam ram_block11a0.clk1_output_clock_enable = "ena1";
defparam ram_block11a0.data_interleave_offset_in_bits = 1;
defparam ram_block11a0.data_interleave_width_in_bits = 1;
defparam ram_block11a0.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a0.operation_mode = "dual_port";
defparam ram_block11a0.port_a_address_clear = "none";
defparam ram_block11a0.port_a_address_width = 8;
defparam ram_block11a0.port_a_data_out_clear = "none";
defparam ram_block11a0.port_a_data_out_clock = "none";
defparam ram_block11a0.port_a_data_width = 1;
defparam ram_block11a0.port_a_first_address = 0;
defparam ram_block11a0.port_a_first_bit_number = 0;
defparam ram_block11a0.port_a_last_address = 255;
defparam ram_block11a0.port_a_logical_ram_depth = 256;
defparam ram_block11a0.port_a_logical_ram_width = 32;
defparam ram_block11a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a0.port_b_address_clear = "clear1";
defparam ram_block11a0.port_b_address_clock = "clock1";
defparam ram_block11a0.port_b_address_width = 8;
defparam ram_block11a0.port_b_data_out_clear = "clear1";
defparam ram_block11a0.port_b_data_out_clock = "clock1";
defparam ram_block11a0.port_b_data_width = 1;
defparam ram_block11a0.port_b_first_address = 0;
defparam ram_block11a0.port_b_first_bit_number = 0;
defparam ram_block11a0.port_b_last_address = 255;
defparam ram_block11a0.port_b_logical_ram_depth = 256;
defparam ram_block11a0.port_b_logical_ram_width = 32;
defparam ram_block11a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a0.port_b_read_enable_clock = "clock1";
defparam ram_block11a0.ram_block_type = "auto";

cyclonev_ram_block ram_block11a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a1.clk0_core_clock_enable = "ena0";
defparam ram_block11a1.clk1_output_clock_enable = "ena1";
defparam ram_block11a1.data_interleave_offset_in_bits = 1;
defparam ram_block11a1.data_interleave_width_in_bits = 1;
defparam ram_block11a1.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a1.operation_mode = "dual_port";
defparam ram_block11a1.port_a_address_clear = "none";
defparam ram_block11a1.port_a_address_width = 8;
defparam ram_block11a1.port_a_data_out_clear = "none";
defparam ram_block11a1.port_a_data_out_clock = "none";
defparam ram_block11a1.port_a_data_width = 1;
defparam ram_block11a1.port_a_first_address = 0;
defparam ram_block11a1.port_a_first_bit_number = 1;
defparam ram_block11a1.port_a_last_address = 255;
defparam ram_block11a1.port_a_logical_ram_depth = 256;
defparam ram_block11a1.port_a_logical_ram_width = 32;
defparam ram_block11a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a1.port_b_address_clear = "clear1";
defparam ram_block11a1.port_b_address_clock = "clock1";
defparam ram_block11a1.port_b_address_width = 8;
defparam ram_block11a1.port_b_data_out_clear = "clear1";
defparam ram_block11a1.port_b_data_out_clock = "clock1";
defparam ram_block11a1.port_b_data_width = 1;
defparam ram_block11a1.port_b_first_address = 0;
defparam ram_block11a1.port_b_first_bit_number = 1;
defparam ram_block11a1.port_b_last_address = 255;
defparam ram_block11a1.port_b_logical_ram_depth = 256;
defparam ram_block11a1.port_b_logical_ram_width = 32;
defparam ram_block11a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a1.port_b_read_enable_clock = "clock1";
defparam ram_block11a1.ram_block_type = "auto";

cyclonev_ram_block ram_block11a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a2.clk0_core_clock_enable = "ena0";
defparam ram_block11a2.clk1_output_clock_enable = "ena1";
defparam ram_block11a2.data_interleave_offset_in_bits = 1;
defparam ram_block11a2.data_interleave_width_in_bits = 1;
defparam ram_block11a2.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a2.operation_mode = "dual_port";
defparam ram_block11a2.port_a_address_clear = "none";
defparam ram_block11a2.port_a_address_width = 8;
defparam ram_block11a2.port_a_data_out_clear = "none";
defparam ram_block11a2.port_a_data_out_clock = "none";
defparam ram_block11a2.port_a_data_width = 1;
defparam ram_block11a2.port_a_first_address = 0;
defparam ram_block11a2.port_a_first_bit_number = 2;
defparam ram_block11a2.port_a_last_address = 255;
defparam ram_block11a2.port_a_logical_ram_depth = 256;
defparam ram_block11a2.port_a_logical_ram_width = 32;
defparam ram_block11a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a2.port_b_address_clear = "clear1";
defparam ram_block11a2.port_b_address_clock = "clock1";
defparam ram_block11a2.port_b_address_width = 8;
defparam ram_block11a2.port_b_data_out_clear = "clear1";
defparam ram_block11a2.port_b_data_out_clock = "clock1";
defparam ram_block11a2.port_b_data_width = 1;
defparam ram_block11a2.port_b_first_address = 0;
defparam ram_block11a2.port_b_first_bit_number = 2;
defparam ram_block11a2.port_b_last_address = 255;
defparam ram_block11a2.port_b_logical_ram_depth = 256;
defparam ram_block11a2.port_b_logical_ram_width = 32;
defparam ram_block11a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a2.port_b_read_enable_clock = "clock1";
defparam ram_block11a2.ram_block_type = "auto";

cyclonev_ram_block ram_block11a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a3.clk0_core_clock_enable = "ena0";
defparam ram_block11a3.clk1_output_clock_enable = "ena1";
defparam ram_block11a3.data_interleave_offset_in_bits = 1;
defparam ram_block11a3.data_interleave_width_in_bits = 1;
defparam ram_block11a3.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a3.operation_mode = "dual_port";
defparam ram_block11a3.port_a_address_clear = "none";
defparam ram_block11a3.port_a_address_width = 8;
defparam ram_block11a3.port_a_data_out_clear = "none";
defparam ram_block11a3.port_a_data_out_clock = "none";
defparam ram_block11a3.port_a_data_width = 1;
defparam ram_block11a3.port_a_first_address = 0;
defparam ram_block11a3.port_a_first_bit_number = 3;
defparam ram_block11a3.port_a_last_address = 255;
defparam ram_block11a3.port_a_logical_ram_depth = 256;
defparam ram_block11a3.port_a_logical_ram_width = 32;
defparam ram_block11a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a3.port_b_address_clear = "clear1";
defparam ram_block11a3.port_b_address_clock = "clock1";
defparam ram_block11a3.port_b_address_width = 8;
defparam ram_block11a3.port_b_data_out_clear = "clear1";
defparam ram_block11a3.port_b_data_out_clock = "clock1";
defparam ram_block11a3.port_b_data_width = 1;
defparam ram_block11a3.port_b_first_address = 0;
defparam ram_block11a3.port_b_first_bit_number = 3;
defparam ram_block11a3.port_b_last_address = 255;
defparam ram_block11a3.port_b_logical_ram_depth = 256;
defparam ram_block11a3.port_b_logical_ram_width = 32;
defparam ram_block11a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a3.port_b_read_enable_clock = "clock1";
defparam ram_block11a3.ram_block_type = "auto";

cyclonev_ram_block ram_block11a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a4.clk0_core_clock_enable = "ena0";
defparam ram_block11a4.clk1_output_clock_enable = "ena1";
defparam ram_block11a4.data_interleave_offset_in_bits = 1;
defparam ram_block11a4.data_interleave_width_in_bits = 1;
defparam ram_block11a4.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a4.operation_mode = "dual_port";
defparam ram_block11a4.port_a_address_clear = "none";
defparam ram_block11a4.port_a_address_width = 8;
defparam ram_block11a4.port_a_data_out_clear = "none";
defparam ram_block11a4.port_a_data_out_clock = "none";
defparam ram_block11a4.port_a_data_width = 1;
defparam ram_block11a4.port_a_first_address = 0;
defparam ram_block11a4.port_a_first_bit_number = 4;
defparam ram_block11a4.port_a_last_address = 255;
defparam ram_block11a4.port_a_logical_ram_depth = 256;
defparam ram_block11a4.port_a_logical_ram_width = 32;
defparam ram_block11a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a4.port_b_address_clear = "clear1";
defparam ram_block11a4.port_b_address_clock = "clock1";
defparam ram_block11a4.port_b_address_width = 8;
defparam ram_block11a4.port_b_data_out_clear = "clear1";
defparam ram_block11a4.port_b_data_out_clock = "clock1";
defparam ram_block11a4.port_b_data_width = 1;
defparam ram_block11a4.port_b_first_address = 0;
defparam ram_block11a4.port_b_first_bit_number = 4;
defparam ram_block11a4.port_b_last_address = 255;
defparam ram_block11a4.port_b_logical_ram_depth = 256;
defparam ram_block11a4.port_b_logical_ram_width = 32;
defparam ram_block11a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a4.port_b_read_enable_clock = "clock1";
defparam ram_block11a4.ram_block_type = "auto";

cyclonev_ram_block ram_block11a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a5.clk0_core_clock_enable = "ena0";
defparam ram_block11a5.clk1_output_clock_enable = "ena1";
defparam ram_block11a5.data_interleave_offset_in_bits = 1;
defparam ram_block11a5.data_interleave_width_in_bits = 1;
defparam ram_block11a5.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a5.operation_mode = "dual_port";
defparam ram_block11a5.port_a_address_clear = "none";
defparam ram_block11a5.port_a_address_width = 8;
defparam ram_block11a5.port_a_data_out_clear = "none";
defparam ram_block11a5.port_a_data_out_clock = "none";
defparam ram_block11a5.port_a_data_width = 1;
defparam ram_block11a5.port_a_first_address = 0;
defparam ram_block11a5.port_a_first_bit_number = 5;
defparam ram_block11a5.port_a_last_address = 255;
defparam ram_block11a5.port_a_logical_ram_depth = 256;
defparam ram_block11a5.port_a_logical_ram_width = 32;
defparam ram_block11a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a5.port_b_address_clear = "clear1";
defparam ram_block11a5.port_b_address_clock = "clock1";
defparam ram_block11a5.port_b_address_width = 8;
defparam ram_block11a5.port_b_data_out_clear = "clear1";
defparam ram_block11a5.port_b_data_out_clock = "clock1";
defparam ram_block11a5.port_b_data_width = 1;
defparam ram_block11a5.port_b_first_address = 0;
defparam ram_block11a5.port_b_first_bit_number = 5;
defparam ram_block11a5.port_b_last_address = 255;
defparam ram_block11a5.port_b_logical_ram_depth = 256;
defparam ram_block11a5.port_b_logical_ram_width = 32;
defparam ram_block11a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a5.port_b_read_enable_clock = "clock1";
defparam ram_block11a5.ram_block_type = "auto";

cyclonev_ram_block ram_block11a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a6.clk0_core_clock_enable = "ena0";
defparam ram_block11a6.clk1_output_clock_enable = "ena1";
defparam ram_block11a6.data_interleave_offset_in_bits = 1;
defparam ram_block11a6.data_interleave_width_in_bits = 1;
defparam ram_block11a6.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a6.operation_mode = "dual_port";
defparam ram_block11a6.port_a_address_clear = "none";
defparam ram_block11a6.port_a_address_width = 8;
defparam ram_block11a6.port_a_data_out_clear = "none";
defparam ram_block11a6.port_a_data_out_clock = "none";
defparam ram_block11a6.port_a_data_width = 1;
defparam ram_block11a6.port_a_first_address = 0;
defparam ram_block11a6.port_a_first_bit_number = 6;
defparam ram_block11a6.port_a_last_address = 255;
defparam ram_block11a6.port_a_logical_ram_depth = 256;
defparam ram_block11a6.port_a_logical_ram_width = 32;
defparam ram_block11a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a6.port_b_address_clear = "clear1";
defparam ram_block11a6.port_b_address_clock = "clock1";
defparam ram_block11a6.port_b_address_width = 8;
defparam ram_block11a6.port_b_data_out_clear = "clear1";
defparam ram_block11a6.port_b_data_out_clock = "clock1";
defparam ram_block11a6.port_b_data_width = 1;
defparam ram_block11a6.port_b_first_address = 0;
defparam ram_block11a6.port_b_first_bit_number = 6;
defparam ram_block11a6.port_b_last_address = 255;
defparam ram_block11a6.port_b_logical_ram_depth = 256;
defparam ram_block11a6.port_b_logical_ram_width = 32;
defparam ram_block11a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a6.port_b_read_enable_clock = "clock1";
defparam ram_block11a6.ram_block_type = "auto";

cyclonev_ram_block ram_block11a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a7.clk0_core_clock_enable = "ena0";
defparam ram_block11a7.clk1_output_clock_enable = "ena1";
defparam ram_block11a7.data_interleave_offset_in_bits = 1;
defparam ram_block11a7.data_interleave_width_in_bits = 1;
defparam ram_block11a7.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a7.operation_mode = "dual_port";
defparam ram_block11a7.port_a_address_clear = "none";
defparam ram_block11a7.port_a_address_width = 8;
defparam ram_block11a7.port_a_data_out_clear = "none";
defparam ram_block11a7.port_a_data_out_clock = "none";
defparam ram_block11a7.port_a_data_width = 1;
defparam ram_block11a7.port_a_first_address = 0;
defparam ram_block11a7.port_a_first_bit_number = 7;
defparam ram_block11a7.port_a_last_address = 255;
defparam ram_block11a7.port_a_logical_ram_depth = 256;
defparam ram_block11a7.port_a_logical_ram_width = 32;
defparam ram_block11a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a7.port_b_address_clear = "clear1";
defparam ram_block11a7.port_b_address_clock = "clock1";
defparam ram_block11a7.port_b_address_width = 8;
defparam ram_block11a7.port_b_data_out_clear = "clear1";
defparam ram_block11a7.port_b_data_out_clock = "clock1";
defparam ram_block11a7.port_b_data_width = 1;
defparam ram_block11a7.port_b_first_address = 0;
defparam ram_block11a7.port_b_first_bit_number = 7;
defparam ram_block11a7.port_b_last_address = 255;
defparam ram_block11a7.port_b_logical_ram_depth = 256;
defparam ram_block11a7.port_b_logical_ram_width = 32;
defparam ram_block11a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a7.port_b_read_enable_clock = "clock1";
defparam ram_block11a7.ram_block_type = "auto";

cyclonev_ram_block ram_block11a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a8.clk0_core_clock_enable = "ena0";
defparam ram_block11a8.clk1_output_clock_enable = "ena1";
defparam ram_block11a8.data_interleave_offset_in_bits = 1;
defparam ram_block11a8.data_interleave_width_in_bits = 1;
defparam ram_block11a8.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a8.operation_mode = "dual_port";
defparam ram_block11a8.port_a_address_clear = "none";
defparam ram_block11a8.port_a_address_width = 8;
defparam ram_block11a8.port_a_data_out_clear = "none";
defparam ram_block11a8.port_a_data_out_clock = "none";
defparam ram_block11a8.port_a_data_width = 1;
defparam ram_block11a8.port_a_first_address = 0;
defparam ram_block11a8.port_a_first_bit_number = 8;
defparam ram_block11a8.port_a_last_address = 255;
defparam ram_block11a8.port_a_logical_ram_depth = 256;
defparam ram_block11a8.port_a_logical_ram_width = 32;
defparam ram_block11a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a8.port_b_address_clear = "clear1";
defparam ram_block11a8.port_b_address_clock = "clock1";
defparam ram_block11a8.port_b_address_width = 8;
defparam ram_block11a8.port_b_data_out_clear = "clear1";
defparam ram_block11a8.port_b_data_out_clock = "clock1";
defparam ram_block11a8.port_b_data_width = 1;
defparam ram_block11a8.port_b_first_address = 0;
defparam ram_block11a8.port_b_first_bit_number = 8;
defparam ram_block11a8.port_b_last_address = 255;
defparam ram_block11a8.port_b_logical_ram_depth = 256;
defparam ram_block11a8.port_b_logical_ram_width = 32;
defparam ram_block11a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a8.port_b_read_enable_clock = "clock1";
defparam ram_block11a8.ram_block_type = "auto";

cyclonev_ram_block ram_block11a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a9.clk0_core_clock_enable = "ena0";
defparam ram_block11a9.clk1_output_clock_enable = "ena1";
defparam ram_block11a9.data_interleave_offset_in_bits = 1;
defparam ram_block11a9.data_interleave_width_in_bits = 1;
defparam ram_block11a9.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a9.operation_mode = "dual_port";
defparam ram_block11a9.port_a_address_clear = "none";
defparam ram_block11a9.port_a_address_width = 8;
defparam ram_block11a9.port_a_data_out_clear = "none";
defparam ram_block11a9.port_a_data_out_clock = "none";
defparam ram_block11a9.port_a_data_width = 1;
defparam ram_block11a9.port_a_first_address = 0;
defparam ram_block11a9.port_a_first_bit_number = 9;
defparam ram_block11a9.port_a_last_address = 255;
defparam ram_block11a9.port_a_logical_ram_depth = 256;
defparam ram_block11a9.port_a_logical_ram_width = 32;
defparam ram_block11a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a9.port_b_address_clear = "clear1";
defparam ram_block11a9.port_b_address_clock = "clock1";
defparam ram_block11a9.port_b_address_width = 8;
defparam ram_block11a9.port_b_data_out_clear = "clear1";
defparam ram_block11a9.port_b_data_out_clock = "clock1";
defparam ram_block11a9.port_b_data_width = 1;
defparam ram_block11a9.port_b_first_address = 0;
defparam ram_block11a9.port_b_first_bit_number = 9;
defparam ram_block11a9.port_b_last_address = 255;
defparam ram_block11a9.port_b_logical_ram_depth = 256;
defparam ram_block11a9.port_b_logical_ram_width = 32;
defparam ram_block11a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a9.port_b_read_enable_clock = "clock1";
defparam ram_block11a9.ram_block_type = "auto";

cyclonev_ram_block ram_block11a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a10.clk0_core_clock_enable = "ena0";
defparam ram_block11a10.clk1_output_clock_enable = "ena1";
defparam ram_block11a10.data_interleave_offset_in_bits = 1;
defparam ram_block11a10.data_interleave_width_in_bits = 1;
defparam ram_block11a10.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a10.operation_mode = "dual_port";
defparam ram_block11a10.port_a_address_clear = "none";
defparam ram_block11a10.port_a_address_width = 8;
defparam ram_block11a10.port_a_data_out_clear = "none";
defparam ram_block11a10.port_a_data_out_clock = "none";
defparam ram_block11a10.port_a_data_width = 1;
defparam ram_block11a10.port_a_first_address = 0;
defparam ram_block11a10.port_a_first_bit_number = 10;
defparam ram_block11a10.port_a_last_address = 255;
defparam ram_block11a10.port_a_logical_ram_depth = 256;
defparam ram_block11a10.port_a_logical_ram_width = 32;
defparam ram_block11a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a10.port_b_address_clear = "clear1";
defparam ram_block11a10.port_b_address_clock = "clock1";
defparam ram_block11a10.port_b_address_width = 8;
defparam ram_block11a10.port_b_data_out_clear = "clear1";
defparam ram_block11a10.port_b_data_out_clock = "clock1";
defparam ram_block11a10.port_b_data_width = 1;
defparam ram_block11a10.port_b_first_address = 0;
defparam ram_block11a10.port_b_first_bit_number = 10;
defparam ram_block11a10.port_b_last_address = 255;
defparam ram_block11a10.port_b_logical_ram_depth = 256;
defparam ram_block11a10.port_b_logical_ram_width = 32;
defparam ram_block11a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a10.port_b_read_enable_clock = "clock1";
defparam ram_block11a10.ram_block_type = "auto";

cyclonev_ram_block ram_block11a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a11.clk0_core_clock_enable = "ena0";
defparam ram_block11a11.clk1_output_clock_enable = "ena1";
defparam ram_block11a11.data_interleave_offset_in_bits = 1;
defparam ram_block11a11.data_interleave_width_in_bits = 1;
defparam ram_block11a11.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a11.operation_mode = "dual_port";
defparam ram_block11a11.port_a_address_clear = "none";
defparam ram_block11a11.port_a_address_width = 8;
defparam ram_block11a11.port_a_data_out_clear = "none";
defparam ram_block11a11.port_a_data_out_clock = "none";
defparam ram_block11a11.port_a_data_width = 1;
defparam ram_block11a11.port_a_first_address = 0;
defparam ram_block11a11.port_a_first_bit_number = 11;
defparam ram_block11a11.port_a_last_address = 255;
defparam ram_block11a11.port_a_logical_ram_depth = 256;
defparam ram_block11a11.port_a_logical_ram_width = 32;
defparam ram_block11a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a11.port_b_address_clear = "clear1";
defparam ram_block11a11.port_b_address_clock = "clock1";
defparam ram_block11a11.port_b_address_width = 8;
defparam ram_block11a11.port_b_data_out_clear = "clear1";
defparam ram_block11a11.port_b_data_out_clock = "clock1";
defparam ram_block11a11.port_b_data_width = 1;
defparam ram_block11a11.port_b_first_address = 0;
defparam ram_block11a11.port_b_first_bit_number = 11;
defparam ram_block11a11.port_b_last_address = 255;
defparam ram_block11a11.port_b_logical_ram_depth = 256;
defparam ram_block11a11.port_b_logical_ram_width = 32;
defparam ram_block11a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a11.port_b_read_enable_clock = "clock1";
defparam ram_block11a11.ram_block_type = "auto";

cyclonev_ram_block ram_block11a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a12.clk0_core_clock_enable = "ena0";
defparam ram_block11a12.clk1_output_clock_enable = "ena1";
defparam ram_block11a12.data_interleave_offset_in_bits = 1;
defparam ram_block11a12.data_interleave_width_in_bits = 1;
defparam ram_block11a12.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a12.operation_mode = "dual_port";
defparam ram_block11a12.port_a_address_clear = "none";
defparam ram_block11a12.port_a_address_width = 8;
defparam ram_block11a12.port_a_data_out_clear = "none";
defparam ram_block11a12.port_a_data_out_clock = "none";
defparam ram_block11a12.port_a_data_width = 1;
defparam ram_block11a12.port_a_first_address = 0;
defparam ram_block11a12.port_a_first_bit_number = 12;
defparam ram_block11a12.port_a_last_address = 255;
defparam ram_block11a12.port_a_logical_ram_depth = 256;
defparam ram_block11a12.port_a_logical_ram_width = 32;
defparam ram_block11a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a12.port_b_address_clear = "clear1";
defparam ram_block11a12.port_b_address_clock = "clock1";
defparam ram_block11a12.port_b_address_width = 8;
defparam ram_block11a12.port_b_data_out_clear = "clear1";
defparam ram_block11a12.port_b_data_out_clock = "clock1";
defparam ram_block11a12.port_b_data_width = 1;
defparam ram_block11a12.port_b_first_address = 0;
defparam ram_block11a12.port_b_first_bit_number = 12;
defparam ram_block11a12.port_b_last_address = 255;
defparam ram_block11a12.port_b_logical_ram_depth = 256;
defparam ram_block11a12.port_b_logical_ram_width = 32;
defparam ram_block11a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a12.port_b_read_enable_clock = "clock1";
defparam ram_block11a12.ram_block_type = "auto";

cyclonev_ram_block ram_block11a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a13.clk0_core_clock_enable = "ena0";
defparam ram_block11a13.clk1_output_clock_enable = "ena1";
defparam ram_block11a13.data_interleave_offset_in_bits = 1;
defparam ram_block11a13.data_interleave_width_in_bits = 1;
defparam ram_block11a13.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a13.operation_mode = "dual_port";
defparam ram_block11a13.port_a_address_clear = "none";
defparam ram_block11a13.port_a_address_width = 8;
defparam ram_block11a13.port_a_data_out_clear = "none";
defparam ram_block11a13.port_a_data_out_clock = "none";
defparam ram_block11a13.port_a_data_width = 1;
defparam ram_block11a13.port_a_first_address = 0;
defparam ram_block11a13.port_a_first_bit_number = 13;
defparam ram_block11a13.port_a_last_address = 255;
defparam ram_block11a13.port_a_logical_ram_depth = 256;
defparam ram_block11a13.port_a_logical_ram_width = 32;
defparam ram_block11a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a13.port_b_address_clear = "clear1";
defparam ram_block11a13.port_b_address_clock = "clock1";
defparam ram_block11a13.port_b_address_width = 8;
defparam ram_block11a13.port_b_data_out_clear = "clear1";
defparam ram_block11a13.port_b_data_out_clock = "clock1";
defparam ram_block11a13.port_b_data_width = 1;
defparam ram_block11a13.port_b_first_address = 0;
defparam ram_block11a13.port_b_first_bit_number = 13;
defparam ram_block11a13.port_b_last_address = 255;
defparam ram_block11a13.port_b_logical_ram_depth = 256;
defparam ram_block11a13.port_b_logical_ram_width = 32;
defparam ram_block11a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a13.port_b_read_enable_clock = "clock1";
defparam ram_block11a13.ram_block_type = "auto";

cyclonev_ram_block ram_block11a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a14.clk0_core_clock_enable = "ena0";
defparam ram_block11a14.clk1_output_clock_enable = "ena1";
defparam ram_block11a14.data_interleave_offset_in_bits = 1;
defparam ram_block11a14.data_interleave_width_in_bits = 1;
defparam ram_block11a14.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a14.operation_mode = "dual_port";
defparam ram_block11a14.port_a_address_clear = "none";
defparam ram_block11a14.port_a_address_width = 8;
defparam ram_block11a14.port_a_data_out_clear = "none";
defparam ram_block11a14.port_a_data_out_clock = "none";
defparam ram_block11a14.port_a_data_width = 1;
defparam ram_block11a14.port_a_first_address = 0;
defparam ram_block11a14.port_a_first_bit_number = 14;
defparam ram_block11a14.port_a_last_address = 255;
defparam ram_block11a14.port_a_logical_ram_depth = 256;
defparam ram_block11a14.port_a_logical_ram_width = 32;
defparam ram_block11a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a14.port_b_address_clear = "clear1";
defparam ram_block11a14.port_b_address_clock = "clock1";
defparam ram_block11a14.port_b_address_width = 8;
defparam ram_block11a14.port_b_data_out_clear = "clear1";
defparam ram_block11a14.port_b_data_out_clock = "clock1";
defparam ram_block11a14.port_b_data_width = 1;
defparam ram_block11a14.port_b_first_address = 0;
defparam ram_block11a14.port_b_first_bit_number = 14;
defparam ram_block11a14.port_b_last_address = 255;
defparam ram_block11a14.port_b_logical_ram_depth = 256;
defparam ram_block11a14.port_b_logical_ram_width = 32;
defparam ram_block11a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a14.port_b_read_enable_clock = "clock1";
defparam ram_block11a14.ram_block_type = "auto";

cyclonev_ram_block ram_block11a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a15.clk0_core_clock_enable = "ena0";
defparam ram_block11a15.clk1_output_clock_enable = "ena1";
defparam ram_block11a15.data_interleave_offset_in_bits = 1;
defparam ram_block11a15.data_interleave_width_in_bits = 1;
defparam ram_block11a15.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a15.operation_mode = "dual_port";
defparam ram_block11a15.port_a_address_clear = "none";
defparam ram_block11a15.port_a_address_width = 8;
defparam ram_block11a15.port_a_data_out_clear = "none";
defparam ram_block11a15.port_a_data_out_clock = "none";
defparam ram_block11a15.port_a_data_width = 1;
defparam ram_block11a15.port_a_first_address = 0;
defparam ram_block11a15.port_a_first_bit_number = 15;
defparam ram_block11a15.port_a_last_address = 255;
defparam ram_block11a15.port_a_logical_ram_depth = 256;
defparam ram_block11a15.port_a_logical_ram_width = 32;
defparam ram_block11a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a15.port_b_address_clear = "clear1";
defparam ram_block11a15.port_b_address_clock = "clock1";
defparam ram_block11a15.port_b_address_width = 8;
defparam ram_block11a15.port_b_data_out_clear = "clear1";
defparam ram_block11a15.port_b_data_out_clock = "clock1";
defparam ram_block11a15.port_b_data_width = 1;
defparam ram_block11a15.port_b_first_address = 0;
defparam ram_block11a15.port_b_first_bit_number = 15;
defparam ram_block11a15.port_b_last_address = 255;
defparam ram_block11a15.port_b_logical_ram_depth = 256;
defparam ram_block11a15.port_b_logical_ram_width = 32;
defparam ram_block11a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a15.port_b_read_enable_clock = "clock1";
defparam ram_block11a15.ram_block_type = "auto";

cyclonev_ram_block ram_block11a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a16.clk0_core_clock_enable = "ena0";
defparam ram_block11a16.clk1_output_clock_enable = "ena1";
defparam ram_block11a16.data_interleave_offset_in_bits = 1;
defparam ram_block11a16.data_interleave_width_in_bits = 1;
defparam ram_block11a16.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a16.operation_mode = "dual_port";
defparam ram_block11a16.port_a_address_clear = "none";
defparam ram_block11a16.port_a_address_width = 8;
defparam ram_block11a16.port_a_data_out_clear = "none";
defparam ram_block11a16.port_a_data_out_clock = "none";
defparam ram_block11a16.port_a_data_width = 1;
defparam ram_block11a16.port_a_first_address = 0;
defparam ram_block11a16.port_a_first_bit_number = 16;
defparam ram_block11a16.port_a_last_address = 255;
defparam ram_block11a16.port_a_logical_ram_depth = 256;
defparam ram_block11a16.port_a_logical_ram_width = 32;
defparam ram_block11a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a16.port_b_address_clear = "clear1";
defparam ram_block11a16.port_b_address_clock = "clock1";
defparam ram_block11a16.port_b_address_width = 8;
defparam ram_block11a16.port_b_data_out_clear = "clear1";
defparam ram_block11a16.port_b_data_out_clock = "clock1";
defparam ram_block11a16.port_b_data_width = 1;
defparam ram_block11a16.port_b_first_address = 0;
defparam ram_block11a16.port_b_first_bit_number = 16;
defparam ram_block11a16.port_b_last_address = 255;
defparam ram_block11a16.port_b_logical_ram_depth = 256;
defparam ram_block11a16.port_b_logical_ram_width = 32;
defparam ram_block11a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a16.port_b_read_enable_clock = "clock1";
defparam ram_block11a16.ram_block_type = "auto";

cyclonev_ram_block ram_block11a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a17.clk0_core_clock_enable = "ena0";
defparam ram_block11a17.clk1_output_clock_enable = "ena1";
defparam ram_block11a17.data_interleave_offset_in_bits = 1;
defparam ram_block11a17.data_interleave_width_in_bits = 1;
defparam ram_block11a17.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a17.operation_mode = "dual_port";
defparam ram_block11a17.port_a_address_clear = "none";
defparam ram_block11a17.port_a_address_width = 8;
defparam ram_block11a17.port_a_data_out_clear = "none";
defparam ram_block11a17.port_a_data_out_clock = "none";
defparam ram_block11a17.port_a_data_width = 1;
defparam ram_block11a17.port_a_first_address = 0;
defparam ram_block11a17.port_a_first_bit_number = 17;
defparam ram_block11a17.port_a_last_address = 255;
defparam ram_block11a17.port_a_logical_ram_depth = 256;
defparam ram_block11a17.port_a_logical_ram_width = 32;
defparam ram_block11a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a17.port_b_address_clear = "clear1";
defparam ram_block11a17.port_b_address_clock = "clock1";
defparam ram_block11a17.port_b_address_width = 8;
defparam ram_block11a17.port_b_data_out_clear = "clear1";
defparam ram_block11a17.port_b_data_out_clock = "clock1";
defparam ram_block11a17.port_b_data_width = 1;
defparam ram_block11a17.port_b_first_address = 0;
defparam ram_block11a17.port_b_first_bit_number = 17;
defparam ram_block11a17.port_b_last_address = 255;
defparam ram_block11a17.port_b_logical_ram_depth = 256;
defparam ram_block11a17.port_b_logical_ram_width = 32;
defparam ram_block11a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a17.port_b_read_enable_clock = "clock1";
defparam ram_block11a17.ram_block_type = "auto";

cyclonev_ram_block ram_block11a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a18.clk0_core_clock_enable = "ena0";
defparam ram_block11a18.clk1_output_clock_enable = "ena1";
defparam ram_block11a18.data_interleave_offset_in_bits = 1;
defparam ram_block11a18.data_interleave_width_in_bits = 1;
defparam ram_block11a18.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a18.operation_mode = "dual_port";
defparam ram_block11a18.port_a_address_clear = "none";
defparam ram_block11a18.port_a_address_width = 8;
defparam ram_block11a18.port_a_data_out_clear = "none";
defparam ram_block11a18.port_a_data_out_clock = "none";
defparam ram_block11a18.port_a_data_width = 1;
defparam ram_block11a18.port_a_first_address = 0;
defparam ram_block11a18.port_a_first_bit_number = 18;
defparam ram_block11a18.port_a_last_address = 255;
defparam ram_block11a18.port_a_logical_ram_depth = 256;
defparam ram_block11a18.port_a_logical_ram_width = 32;
defparam ram_block11a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a18.port_b_address_clear = "clear1";
defparam ram_block11a18.port_b_address_clock = "clock1";
defparam ram_block11a18.port_b_address_width = 8;
defparam ram_block11a18.port_b_data_out_clear = "clear1";
defparam ram_block11a18.port_b_data_out_clock = "clock1";
defparam ram_block11a18.port_b_data_width = 1;
defparam ram_block11a18.port_b_first_address = 0;
defparam ram_block11a18.port_b_first_bit_number = 18;
defparam ram_block11a18.port_b_last_address = 255;
defparam ram_block11a18.port_b_logical_ram_depth = 256;
defparam ram_block11a18.port_b_logical_ram_width = 32;
defparam ram_block11a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a18.port_b_read_enable_clock = "clock1";
defparam ram_block11a18.ram_block_type = "auto";

cyclonev_ram_block ram_block11a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a19.clk0_core_clock_enable = "ena0";
defparam ram_block11a19.clk1_output_clock_enable = "ena1";
defparam ram_block11a19.data_interleave_offset_in_bits = 1;
defparam ram_block11a19.data_interleave_width_in_bits = 1;
defparam ram_block11a19.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a19.operation_mode = "dual_port";
defparam ram_block11a19.port_a_address_clear = "none";
defparam ram_block11a19.port_a_address_width = 8;
defparam ram_block11a19.port_a_data_out_clear = "none";
defparam ram_block11a19.port_a_data_out_clock = "none";
defparam ram_block11a19.port_a_data_width = 1;
defparam ram_block11a19.port_a_first_address = 0;
defparam ram_block11a19.port_a_first_bit_number = 19;
defparam ram_block11a19.port_a_last_address = 255;
defparam ram_block11a19.port_a_logical_ram_depth = 256;
defparam ram_block11a19.port_a_logical_ram_width = 32;
defparam ram_block11a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a19.port_b_address_clear = "clear1";
defparam ram_block11a19.port_b_address_clock = "clock1";
defparam ram_block11a19.port_b_address_width = 8;
defparam ram_block11a19.port_b_data_out_clear = "clear1";
defparam ram_block11a19.port_b_data_out_clock = "clock1";
defparam ram_block11a19.port_b_data_width = 1;
defparam ram_block11a19.port_b_first_address = 0;
defparam ram_block11a19.port_b_first_bit_number = 19;
defparam ram_block11a19.port_b_last_address = 255;
defparam ram_block11a19.port_b_logical_ram_depth = 256;
defparam ram_block11a19.port_b_logical_ram_width = 32;
defparam ram_block11a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a19.port_b_read_enable_clock = "clock1";
defparam ram_block11a19.ram_block_type = "auto";

cyclonev_ram_block ram_block11a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a20.clk0_core_clock_enable = "ena0";
defparam ram_block11a20.clk1_output_clock_enable = "ena1";
defparam ram_block11a20.data_interleave_offset_in_bits = 1;
defparam ram_block11a20.data_interleave_width_in_bits = 1;
defparam ram_block11a20.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a20.operation_mode = "dual_port";
defparam ram_block11a20.port_a_address_clear = "none";
defparam ram_block11a20.port_a_address_width = 8;
defparam ram_block11a20.port_a_data_out_clear = "none";
defparam ram_block11a20.port_a_data_out_clock = "none";
defparam ram_block11a20.port_a_data_width = 1;
defparam ram_block11a20.port_a_first_address = 0;
defparam ram_block11a20.port_a_first_bit_number = 20;
defparam ram_block11a20.port_a_last_address = 255;
defparam ram_block11a20.port_a_logical_ram_depth = 256;
defparam ram_block11a20.port_a_logical_ram_width = 32;
defparam ram_block11a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a20.port_b_address_clear = "clear1";
defparam ram_block11a20.port_b_address_clock = "clock1";
defparam ram_block11a20.port_b_address_width = 8;
defparam ram_block11a20.port_b_data_out_clear = "clear1";
defparam ram_block11a20.port_b_data_out_clock = "clock1";
defparam ram_block11a20.port_b_data_width = 1;
defparam ram_block11a20.port_b_first_address = 0;
defparam ram_block11a20.port_b_first_bit_number = 20;
defparam ram_block11a20.port_b_last_address = 255;
defparam ram_block11a20.port_b_logical_ram_depth = 256;
defparam ram_block11a20.port_b_logical_ram_width = 32;
defparam ram_block11a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a20.port_b_read_enable_clock = "clock1";
defparam ram_block11a20.ram_block_type = "auto";

cyclonev_ram_block ram_block11a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a21.clk0_core_clock_enable = "ena0";
defparam ram_block11a21.clk1_output_clock_enable = "ena1";
defparam ram_block11a21.data_interleave_offset_in_bits = 1;
defparam ram_block11a21.data_interleave_width_in_bits = 1;
defparam ram_block11a21.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a21.operation_mode = "dual_port";
defparam ram_block11a21.port_a_address_clear = "none";
defparam ram_block11a21.port_a_address_width = 8;
defparam ram_block11a21.port_a_data_out_clear = "none";
defparam ram_block11a21.port_a_data_out_clock = "none";
defparam ram_block11a21.port_a_data_width = 1;
defparam ram_block11a21.port_a_first_address = 0;
defparam ram_block11a21.port_a_first_bit_number = 21;
defparam ram_block11a21.port_a_last_address = 255;
defparam ram_block11a21.port_a_logical_ram_depth = 256;
defparam ram_block11a21.port_a_logical_ram_width = 32;
defparam ram_block11a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a21.port_b_address_clear = "clear1";
defparam ram_block11a21.port_b_address_clock = "clock1";
defparam ram_block11a21.port_b_address_width = 8;
defparam ram_block11a21.port_b_data_out_clear = "clear1";
defparam ram_block11a21.port_b_data_out_clock = "clock1";
defparam ram_block11a21.port_b_data_width = 1;
defparam ram_block11a21.port_b_first_address = 0;
defparam ram_block11a21.port_b_first_bit_number = 21;
defparam ram_block11a21.port_b_last_address = 255;
defparam ram_block11a21.port_b_logical_ram_depth = 256;
defparam ram_block11a21.port_b_logical_ram_width = 32;
defparam ram_block11a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a21.port_b_read_enable_clock = "clock1";
defparam ram_block11a21.ram_block_type = "auto";

cyclonev_ram_block ram_block11a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a22.clk0_core_clock_enable = "ena0";
defparam ram_block11a22.clk1_output_clock_enable = "ena1";
defparam ram_block11a22.data_interleave_offset_in_bits = 1;
defparam ram_block11a22.data_interleave_width_in_bits = 1;
defparam ram_block11a22.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a22.operation_mode = "dual_port";
defparam ram_block11a22.port_a_address_clear = "none";
defparam ram_block11a22.port_a_address_width = 8;
defparam ram_block11a22.port_a_data_out_clear = "none";
defparam ram_block11a22.port_a_data_out_clock = "none";
defparam ram_block11a22.port_a_data_width = 1;
defparam ram_block11a22.port_a_first_address = 0;
defparam ram_block11a22.port_a_first_bit_number = 22;
defparam ram_block11a22.port_a_last_address = 255;
defparam ram_block11a22.port_a_logical_ram_depth = 256;
defparam ram_block11a22.port_a_logical_ram_width = 32;
defparam ram_block11a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a22.port_b_address_clear = "clear1";
defparam ram_block11a22.port_b_address_clock = "clock1";
defparam ram_block11a22.port_b_address_width = 8;
defparam ram_block11a22.port_b_data_out_clear = "clear1";
defparam ram_block11a22.port_b_data_out_clock = "clock1";
defparam ram_block11a22.port_b_data_width = 1;
defparam ram_block11a22.port_b_first_address = 0;
defparam ram_block11a22.port_b_first_bit_number = 22;
defparam ram_block11a22.port_b_last_address = 255;
defparam ram_block11a22.port_b_logical_ram_depth = 256;
defparam ram_block11a22.port_b_logical_ram_width = 32;
defparam ram_block11a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a22.port_b_read_enable_clock = "clock1";
defparam ram_block11a22.ram_block_type = "auto";

cyclonev_ram_block ram_block11a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a23.clk0_core_clock_enable = "ena0";
defparam ram_block11a23.clk1_output_clock_enable = "ena1";
defparam ram_block11a23.data_interleave_offset_in_bits = 1;
defparam ram_block11a23.data_interleave_width_in_bits = 1;
defparam ram_block11a23.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a23.operation_mode = "dual_port";
defparam ram_block11a23.port_a_address_clear = "none";
defparam ram_block11a23.port_a_address_width = 8;
defparam ram_block11a23.port_a_data_out_clear = "none";
defparam ram_block11a23.port_a_data_out_clock = "none";
defparam ram_block11a23.port_a_data_width = 1;
defparam ram_block11a23.port_a_first_address = 0;
defparam ram_block11a23.port_a_first_bit_number = 23;
defparam ram_block11a23.port_a_last_address = 255;
defparam ram_block11a23.port_a_logical_ram_depth = 256;
defparam ram_block11a23.port_a_logical_ram_width = 32;
defparam ram_block11a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a23.port_b_address_clear = "clear1";
defparam ram_block11a23.port_b_address_clock = "clock1";
defparam ram_block11a23.port_b_address_width = 8;
defparam ram_block11a23.port_b_data_out_clear = "clear1";
defparam ram_block11a23.port_b_data_out_clock = "clock1";
defparam ram_block11a23.port_b_data_width = 1;
defparam ram_block11a23.port_b_first_address = 0;
defparam ram_block11a23.port_b_first_bit_number = 23;
defparam ram_block11a23.port_b_last_address = 255;
defparam ram_block11a23.port_b_logical_ram_depth = 256;
defparam ram_block11a23.port_b_logical_ram_width = 32;
defparam ram_block11a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a23.port_b_read_enable_clock = "clock1";
defparam ram_block11a23.ram_block_type = "auto";

cyclonev_ram_block ram_block11a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a24.clk0_core_clock_enable = "ena0";
defparam ram_block11a24.clk1_output_clock_enable = "ena1";
defparam ram_block11a24.data_interleave_offset_in_bits = 1;
defparam ram_block11a24.data_interleave_width_in_bits = 1;
defparam ram_block11a24.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a24.operation_mode = "dual_port";
defparam ram_block11a24.port_a_address_clear = "none";
defparam ram_block11a24.port_a_address_width = 8;
defparam ram_block11a24.port_a_data_out_clear = "none";
defparam ram_block11a24.port_a_data_out_clock = "none";
defparam ram_block11a24.port_a_data_width = 1;
defparam ram_block11a24.port_a_first_address = 0;
defparam ram_block11a24.port_a_first_bit_number = 24;
defparam ram_block11a24.port_a_last_address = 255;
defparam ram_block11a24.port_a_logical_ram_depth = 256;
defparam ram_block11a24.port_a_logical_ram_width = 32;
defparam ram_block11a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a24.port_b_address_clear = "clear1";
defparam ram_block11a24.port_b_address_clock = "clock1";
defparam ram_block11a24.port_b_address_width = 8;
defparam ram_block11a24.port_b_data_out_clear = "clear1";
defparam ram_block11a24.port_b_data_out_clock = "clock1";
defparam ram_block11a24.port_b_data_width = 1;
defparam ram_block11a24.port_b_first_address = 0;
defparam ram_block11a24.port_b_first_bit_number = 24;
defparam ram_block11a24.port_b_last_address = 255;
defparam ram_block11a24.port_b_logical_ram_depth = 256;
defparam ram_block11a24.port_b_logical_ram_width = 32;
defparam ram_block11a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a24.port_b_read_enable_clock = "clock1";
defparam ram_block11a24.ram_block_type = "auto";

cyclonev_ram_block ram_block11a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a25.clk0_core_clock_enable = "ena0";
defparam ram_block11a25.clk1_output_clock_enable = "ena1";
defparam ram_block11a25.data_interleave_offset_in_bits = 1;
defparam ram_block11a25.data_interleave_width_in_bits = 1;
defparam ram_block11a25.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a25.operation_mode = "dual_port";
defparam ram_block11a25.port_a_address_clear = "none";
defparam ram_block11a25.port_a_address_width = 8;
defparam ram_block11a25.port_a_data_out_clear = "none";
defparam ram_block11a25.port_a_data_out_clock = "none";
defparam ram_block11a25.port_a_data_width = 1;
defparam ram_block11a25.port_a_first_address = 0;
defparam ram_block11a25.port_a_first_bit_number = 25;
defparam ram_block11a25.port_a_last_address = 255;
defparam ram_block11a25.port_a_logical_ram_depth = 256;
defparam ram_block11a25.port_a_logical_ram_width = 32;
defparam ram_block11a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a25.port_b_address_clear = "clear1";
defparam ram_block11a25.port_b_address_clock = "clock1";
defparam ram_block11a25.port_b_address_width = 8;
defparam ram_block11a25.port_b_data_out_clear = "clear1";
defparam ram_block11a25.port_b_data_out_clock = "clock1";
defparam ram_block11a25.port_b_data_width = 1;
defparam ram_block11a25.port_b_first_address = 0;
defparam ram_block11a25.port_b_first_bit_number = 25;
defparam ram_block11a25.port_b_last_address = 255;
defparam ram_block11a25.port_b_logical_ram_depth = 256;
defparam ram_block11a25.port_b_logical_ram_width = 32;
defparam ram_block11a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a25.port_b_read_enable_clock = "clock1";
defparam ram_block11a25.ram_block_type = "auto";

cyclonev_ram_block ram_block11a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a26.clk0_core_clock_enable = "ena0";
defparam ram_block11a26.clk1_output_clock_enable = "ena1";
defparam ram_block11a26.data_interleave_offset_in_bits = 1;
defparam ram_block11a26.data_interleave_width_in_bits = 1;
defparam ram_block11a26.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a26.operation_mode = "dual_port";
defparam ram_block11a26.port_a_address_clear = "none";
defparam ram_block11a26.port_a_address_width = 8;
defparam ram_block11a26.port_a_data_out_clear = "none";
defparam ram_block11a26.port_a_data_out_clock = "none";
defparam ram_block11a26.port_a_data_width = 1;
defparam ram_block11a26.port_a_first_address = 0;
defparam ram_block11a26.port_a_first_bit_number = 26;
defparam ram_block11a26.port_a_last_address = 255;
defparam ram_block11a26.port_a_logical_ram_depth = 256;
defparam ram_block11a26.port_a_logical_ram_width = 32;
defparam ram_block11a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a26.port_b_address_clear = "clear1";
defparam ram_block11a26.port_b_address_clock = "clock1";
defparam ram_block11a26.port_b_address_width = 8;
defparam ram_block11a26.port_b_data_out_clear = "clear1";
defparam ram_block11a26.port_b_data_out_clock = "clock1";
defparam ram_block11a26.port_b_data_width = 1;
defparam ram_block11a26.port_b_first_address = 0;
defparam ram_block11a26.port_b_first_bit_number = 26;
defparam ram_block11a26.port_b_last_address = 255;
defparam ram_block11a26.port_b_logical_ram_depth = 256;
defparam ram_block11a26.port_b_logical_ram_width = 32;
defparam ram_block11a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a26.port_b_read_enable_clock = "clock1";
defparam ram_block11a26.ram_block_type = "auto";

cyclonev_ram_block ram_block11a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a27.clk0_core_clock_enable = "ena0";
defparam ram_block11a27.clk1_output_clock_enable = "ena1";
defparam ram_block11a27.data_interleave_offset_in_bits = 1;
defparam ram_block11a27.data_interleave_width_in_bits = 1;
defparam ram_block11a27.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a27.operation_mode = "dual_port";
defparam ram_block11a27.port_a_address_clear = "none";
defparam ram_block11a27.port_a_address_width = 8;
defparam ram_block11a27.port_a_data_out_clear = "none";
defparam ram_block11a27.port_a_data_out_clock = "none";
defparam ram_block11a27.port_a_data_width = 1;
defparam ram_block11a27.port_a_first_address = 0;
defparam ram_block11a27.port_a_first_bit_number = 27;
defparam ram_block11a27.port_a_last_address = 255;
defparam ram_block11a27.port_a_logical_ram_depth = 256;
defparam ram_block11a27.port_a_logical_ram_width = 32;
defparam ram_block11a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a27.port_b_address_clear = "clear1";
defparam ram_block11a27.port_b_address_clock = "clock1";
defparam ram_block11a27.port_b_address_width = 8;
defparam ram_block11a27.port_b_data_out_clear = "clear1";
defparam ram_block11a27.port_b_data_out_clock = "clock1";
defparam ram_block11a27.port_b_data_width = 1;
defparam ram_block11a27.port_b_first_address = 0;
defparam ram_block11a27.port_b_first_bit_number = 27;
defparam ram_block11a27.port_b_last_address = 255;
defparam ram_block11a27.port_b_logical_ram_depth = 256;
defparam ram_block11a27.port_b_logical_ram_width = 32;
defparam ram_block11a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a27.port_b_read_enable_clock = "clock1";
defparam ram_block11a27.ram_block_type = "auto";

cyclonev_ram_block ram_block11a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a28.clk0_core_clock_enable = "ena0";
defparam ram_block11a28.clk1_output_clock_enable = "ena1";
defparam ram_block11a28.data_interleave_offset_in_bits = 1;
defparam ram_block11a28.data_interleave_width_in_bits = 1;
defparam ram_block11a28.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a28.operation_mode = "dual_port";
defparam ram_block11a28.port_a_address_clear = "none";
defparam ram_block11a28.port_a_address_width = 8;
defparam ram_block11a28.port_a_data_out_clear = "none";
defparam ram_block11a28.port_a_data_out_clock = "none";
defparam ram_block11a28.port_a_data_width = 1;
defparam ram_block11a28.port_a_first_address = 0;
defparam ram_block11a28.port_a_first_bit_number = 28;
defparam ram_block11a28.port_a_last_address = 255;
defparam ram_block11a28.port_a_logical_ram_depth = 256;
defparam ram_block11a28.port_a_logical_ram_width = 32;
defparam ram_block11a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a28.port_b_address_clear = "clear1";
defparam ram_block11a28.port_b_address_clock = "clock1";
defparam ram_block11a28.port_b_address_width = 8;
defparam ram_block11a28.port_b_data_out_clear = "clear1";
defparam ram_block11a28.port_b_data_out_clock = "clock1";
defparam ram_block11a28.port_b_data_width = 1;
defparam ram_block11a28.port_b_first_address = 0;
defparam ram_block11a28.port_b_first_bit_number = 28;
defparam ram_block11a28.port_b_last_address = 255;
defparam ram_block11a28.port_b_logical_ram_depth = 256;
defparam ram_block11a28.port_b_logical_ram_width = 32;
defparam ram_block11a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a28.port_b_read_enable_clock = "clock1";
defparam ram_block11a28.ram_block_type = "auto";

cyclonev_ram_block ram_block11a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a29.clk0_core_clock_enable = "ena0";
defparam ram_block11a29.clk1_output_clock_enable = "ena1";
defparam ram_block11a29.data_interleave_offset_in_bits = 1;
defparam ram_block11a29.data_interleave_width_in_bits = 1;
defparam ram_block11a29.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a29.operation_mode = "dual_port";
defparam ram_block11a29.port_a_address_clear = "none";
defparam ram_block11a29.port_a_address_width = 8;
defparam ram_block11a29.port_a_data_out_clear = "none";
defparam ram_block11a29.port_a_data_out_clock = "none";
defparam ram_block11a29.port_a_data_width = 1;
defparam ram_block11a29.port_a_first_address = 0;
defparam ram_block11a29.port_a_first_bit_number = 29;
defparam ram_block11a29.port_a_last_address = 255;
defparam ram_block11a29.port_a_logical_ram_depth = 256;
defparam ram_block11a29.port_a_logical_ram_width = 32;
defparam ram_block11a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a29.port_b_address_clear = "clear1";
defparam ram_block11a29.port_b_address_clock = "clock1";
defparam ram_block11a29.port_b_address_width = 8;
defparam ram_block11a29.port_b_data_out_clear = "clear1";
defparam ram_block11a29.port_b_data_out_clock = "clock1";
defparam ram_block11a29.port_b_data_width = 1;
defparam ram_block11a29.port_b_first_address = 0;
defparam ram_block11a29.port_b_first_bit_number = 29;
defparam ram_block11a29.port_b_last_address = 255;
defparam ram_block11a29.port_b_logical_ram_depth = 256;
defparam ram_block11a29.port_b_logical_ram_width = 32;
defparam ram_block11a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a29.port_b_read_enable_clock = "clock1";
defparam ram_block11a29.ram_block_type = "auto";

cyclonev_ram_block ram_block11a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a30.clk0_core_clock_enable = "ena0";
defparam ram_block11a30.clk1_output_clock_enable = "ena1";
defparam ram_block11a30.data_interleave_offset_in_bits = 1;
defparam ram_block11a30.data_interleave_width_in_bits = 1;
defparam ram_block11a30.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a30.operation_mode = "dual_port";
defparam ram_block11a30.port_a_address_clear = "none";
defparam ram_block11a30.port_a_address_width = 8;
defparam ram_block11a30.port_a_data_out_clear = "none";
defparam ram_block11a30.port_a_data_out_clock = "none";
defparam ram_block11a30.port_a_data_width = 1;
defparam ram_block11a30.port_a_first_address = 0;
defparam ram_block11a30.port_a_first_bit_number = 30;
defparam ram_block11a30.port_a_last_address = 255;
defparam ram_block11a30.port_a_logical_ram_depth = 256;
defparam ram_block11a30.port_a_logical_ram_width = 32;
defparam ram_block11a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a30.port_b_address_clear = "clear1";
defparam ram_block11a30.port_b_address_clock = "clock1";
defparam ram_block11a30.port_b_address_width = 8;
defparam ram_block11a30.port_b_data_out_clear = "clear1";
defparam ram_block11a30.port_b_data_out_clock = "clock1";
defparam ram_block11a30.port_b_data_width = 1;
defparam ram_block11a30.port_b_first_address = 0;
defparam ram_block11a30.port_b_first_bit_number = 30;
defparam ram_block11a30.port_b_last_address = 255;
defparam ram_block11a30.port_b_logical_ram_depth = 256;
defparam ram_block11a30.port_b_logical_ram_width = 32;
defparam ram_block11a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a30.port_b_read_enable_clock = "clock1";
defparam ram_block11a30.ram_block_type = "auto";

cyclonev_ram_block ram_block11a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(!addressstall_b),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(addressstall_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(!aclr1),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block11a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block11a31.clk0_core_clock_enable = "ena0";
defparam ram_block11a31.clk1_output_clock_enable = "ena1";
defparam ram_block11a31.data_interleave_offset_in_bits = 1;
defparam ram_block11a31.data_interleave_width_in_bits = 1;
defparam ram_block11a31.logical_ram_name = "Computer_System_fifo_HPS_to_FPGA:fifo_hps_to_fpga|Computer_System_fifo_HPS_to_FPGA_dcfifo_with_controls:the_dcfifo_with_controls|Computer_System_fifo_HPS_to_FPGA_dual_clock_fifo:the_dcfifo|dcfifo:dual_clock_fifo|dcfifo_k482:auto_generated|altsyncram_26d1:fifo_ram|ALTSYNCRAM";
defparam ram_block11a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block11a31.operation_mode = "dual_port";
defparam ram_block11a31.port_a_address_clear = "none";
defparam ram_block11a31.port_a_address_width = 8;
defparam ram_block11a31.port_a_data_out_clear = "none";
defparam ram_block11a31.port_a_data_out_clock = "none";
defparam ram_block11a31.port_a_data_width = 1;
defparam ram_block11a31.port_a_first_address = 0;
defparam ram_block11a31.port_a_first_bit_number = 31;
defparam ram_block11a31.port_a_last_address = 255;
defparam ram_block11a31.port_a_logical_ram_depth = 256;
defparam ram_block11a31.port_a_logical_ram_width = 32;
defparam ram_block11a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a31.port_b_address_clear = "clear1";
defparam ram_block11a31.port_b_address_clock = "clock1";
defparam ram_block11a31.port_b_address_width = 8;
defparam ram_block11a31.port_b_data_out_clear = "clear1";
defparam ram_block11a31.port_b_data_out_clock = "clock1";
defparam ram_block11a31.port_b_data_width = 1;
defparam ram_block11a31.port_b_first_address = 0;
defparam ram_block11a31.port_b_first_bit_number = 31;
defparam ram_block11a31.port_b_last_address = 255;
defparam ram_block11a31.port_b_logical_ram_depth = 256;
defparam ram_block11a31.port_b_logical_ram_width = 32;
defparam ram_block11a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block11a31.port_b_read_enable_clock = "clock1";
defparam ram_block11a31.ram_block_type = "auto";

endmodule

module Computer_System_cmpr_1v5 (
	rdptr_g_1,
	dffe17a_1,
	data_wire_2,
	aneb_result_wire_0,
	aneb_result_wire_01,
	rdptr_g_8,
	dffe17a_8,
	rdptr_g_7,
	dffe17a_7,
	aneb_result_wire_02,
	aneb_result_wire_03)/* synthesis synthesis_greybox=0 */;
input 	rdptr_g_1;
input 	dffe17a_1;
output 	data_wire_2;
input 	aneb_result_wire_0;
input 	aneb_result_wire_01;
input 	rdptr_g_8;
input 	dffe17a_8;
input 	rdptr_g_7;
input 	dffe17a_7;
output 	aneb_result_wire_02;
output 	aneb_result_wire_03;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \data_wire[2]~0 (
	.dataa(!rdptr_g_1),
	.datab(!dffe17a_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(data_wire_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_wire[2]~0 .extended_lut = "off";
defparam \data_wire[2]~0 .lut_mask = 64'h6666666666666666;
defparam \data_wire[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \aneb_result_wire[0]~0 (
	.dataa(!rdptr_g_8),
	.datab(!dffe17a_8),
	.datac(!rdptr_g_7),
	.datad(!dffe17a_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(aneb_result_wire_02),
	.sumout(),
	.cout(),
	.shareout());
defparam \aneb_result_wire[0]~0 .extended_lut = "off";
defparam \aneb_result_wire[0]~0 .lut_mask = 64'h9009900990099009;
defparam \aneb_result_wire[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \aneb_result_wire[0] (
	.dataa(!data_wire_2),
	.datab(!aneb_result_wire_0),
	.datac(!aneb_result_wire_01),
	.datad(!aneb_result_wire_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(aneb_result_wire_03),
	.sumout(),
	.cout(),
	.shareout());
defparam \aneb_result_wire[0] .extended_lut = "off";
defparam \aneb_result_wire[0] .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \aneb_result_wire[0] .shared_arith = "off";

endmodule

module Computer_System_cmpr_1v5_1 (
	data_wire_2,
	rdptr_g_6,
	dffe17a_6,
	rdptr_g_4,
	dffe17a_4,
	rdptr_g_5,
	dffe17a_5,
	aneb_result_wire_0,
	rdptr_g_2,
	dffe17a_2,
	rdptr_g_3,
	dffe17a_3,
	rdptr_g_0,
	dffe17a_0,
	aneb_result_wire_01,
	rdptr_g_8,
	dffe17a_8,
	rdptr_g_7,
	dffe17a_7,
	aneb_result_wire_02)/* synthesis synthesis_greybox=0 */;
input 	data_wire_2;
input 	rdptr_g_6;
input 	dffe17a_6;
input 	rdptr_g_4;
input 	dffe17a_4;
input 	rdptr_g_5;
input 	dffe17a_5;
output 	aneb_result_wire_0;
input 	rdptr_g_2;
input 	dffe17a_2;
input 	rdptr_g_3;
input 	dffe17a_3;
input 	rdptr_g_0;
input 	dffe17a_0;
output 	aneb_result_wire_01;
input 	rdptr_g_8;
input 	dffe17a_8;
input 	rdptr_g_7;
input 	dffe17a_7;
output 	aneb_result_wire_02;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \aneb_result_wire[0]~2_combout ;


cyclonev_lcell_comb \aneb_result_wire[0]~0 (
	.dataa(!rdptr_g_6),
	.datab(!dffe17a_6),
	.datac(!rdptr_g_4),
	.datad(!dffe17a_4),
	.datae(!rdptr_g_5),
	.dataf(!dffe17a_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(aneb_result_wire_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \aneb_result_wire[0]~0 .extended_lut = "off";
defparam \aneb_result_wire[0]~0 .lut_mask = 64'h9009000000009009;
defparam \aneb_result_wire[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \aneb_result_wire[0]~1 (
	.dataa(!rdptr_g_2),
	.datab(!dffe17a_2),
	.datac(!rdptr_g_3),
	.datad(!dffe17a_3),
	.datae(!rdptr_g_0),
	.dataf(!dffe17a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(aneb_result_wire_01),
	.sumout(),
	.cout(),
	.shareout());
defparam \aneb_result_wire[0]~1 .extended_lut = "off";
defparam \aneb_result_wire[0]~1 .lut_mask = 64'h9009000000009009;
defparam \aneb_result_wire[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \aneb_result_wire[0]~3 (
	.dataa(!data_wire_2),
	.datab(!aneb_result_wire_0),
	.datac(!aneb_result_wire_01),
	.datad(!\aneb_result_wire[0]~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(aneb_result_wire_02),
	.sumout(),
	.cout(),
	.shareout());
defparam \aneb_result_wire[0]~3 .extended_lut = "off";
defparam \aneb_result_wire[0]~3 .lut_mask = 64'h0002000200020002;
defparam \aneb_result_wire[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \aneb_result_wire[0]~2 (
	.dataa(!rdptr_g_8),
	.datab(!dffe17a_8),
	.datac(!rdptr_g_7),
	.datad(!dffe17a_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aneb_result_wire[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aneb_result_wire[0]~2 .extended_lut = "off";
defparam \aneb_result_wire[0]~2 .lut_mask = 64'h0660066006600660;
defparam \aneb_result_wire[0]~2 .shared_arith = "off";

endmodule

module Computer_System_cmpr_1v5_2 (
	wrptr_g_1,
	dffe20a_1,
	aneb_result_wire_0,
	aneb_result_wire_01,
	wrptr_g_8,
	dffe20a_8,
	wrptr_g_7,
	dffe20a_7,
	aneb_result_wire_02)/* synthesis synthesis_greybox=0 */;
input 	wrptr_g_1;
input 	dffe20a_1;
input 	aneb_result_wire_0;
input 	aneb_result_wire_01;
input 	wrptr_g_8;
input 	dffe20a_8;
input 	wrptr_g_7;
input 	dffe20a_7;
output 	aneb_result_wire_02;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \aneb_result_wire[0]~0_combout ;


cyclonev_lcell_comb \aneb_result_wire[0] (
	.dataa(!wrptr_g_1),
	.datab(!dffe20a_1),
	.datac(!aneb_result_wire_0),
	.datad(!aneb_result_wire_01),
	.datae(!\aneb_result_wire[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(aneb_result_wire_02),
	.sumout(),
	.cout(),
	.shareout());
defparam \aneb_result_wire[0] .extended_lut = "off";
defparam \aneb_result_wire[0] .lut_mask = 64'hFFFFFFF6FFFFFFF6;
defparam \aneb_result_wire[0] .shared_arith = "off";

cyclonev_lcell_comb \aneb_result_wire[0]~0 (
	.dataa(!wrptr_g_8),
	.datab(!dffe20a_8),
	.datac(!wrptr_g_7),
	.datad(!dffe20a_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aneb_result_wire[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aneb_result_wire[0]~0 .extended_lut = "off";
defparam \aneb_result_wire[0]~0 .lut_mask = 64'h9009900990099009;
defparam \aneb_result_wire[0]~0 .shared_arith = "off";

endmodule

module Computer_System_cmpr_1v5_3 (
	wrptr_g_6,
	dffe20a_6,
	wrptr_g_4,
	dffe20a_4,
	wrptr_g_5,
	dffe20a_5,
	aneb_result_wire_0,
	wrptr_g_2,
	dffe20a_2,
	wrptr_g_3,
	dffe20a_3,
	wrptr_g_0,
	dffe20a_0,
	aneb_result_wire_01,
	wrptr_g_8,
	dffe20a_8,
	wrptr_g_7,
	dffe20a_7,
	aneb_result_wire_02)/* synthesis synthesis_greybox=0 */;
input 	wrptr_g_6;
input 	dffe20a_6;
input 	wrptr_g_4;
input 	dffe20a_4;
input 	wrptr_g_5;
input 	dffe20a_5;
output 	aneb_result_wire_0;
input 	wrptr_g_2;
input 	dffe20a_2;
input 	wrptr_g_3;
input 	dffe20a_3;
input 	wrptr_g_0;
input 	dffe20a_0;
output 	aneb_result_wire_01;
input 	wrptr_g_8;
input 	dffe20a_8;
input 	wrptr_g_7;
input 	dffe20a_7;
output 	aneb_result_wire_02;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \aneb_result_wire[0]~0 (
	.dataa(!wrptr_g_6),
	.datab(!dffe20a_6),
	.datac(!wrptr_g_4),
	.datad(!dffe20a_4),
	.datae(!wrptr_g_5),
	.dataf(!dffe20a_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(aneb_result_wire_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \aneb_result_wire[0]~0 .extended_lut = "off";
defparam \aneb_result_wire[0]~0 .lut_mask = 64'h9009000000009009;
defparam \aneb_result_wire[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \aneb_result_wire[0]~1 (
	.dataa(!wrptr_g_2),
	.datab(!dffe20a_2),
	.datac(!wrptr_g_3),
	.datad(!dffe20a_3),
	.datae(!wrptr_g_0),
	.dataf(!dffe20a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(aneb_result_wire_01),
	.sumout(),
	.cout(),
	.shareout());
defparam \aneb_result_wire[0]~1 .extended_lut = "off";
defparam \aneb_result_wire[0]~1 .lut_mask = 64'h9009000000009009;
defparam \aneb_result_wire[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \aneb_result_wire[0]~2 (
	.dataa(!wrptr_g_8),
	.datab(!dffe20a_8),
	.datac(!wrptr_g_7),
	.datad(!dffe20a_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(aneb_result_wire_02),
	.sumout(),
	.cout(),
	.shareout());
defparam \aneb_result_wire[0]~2 .extended_lut = "off";
defparam \aneb_result_wire[0]~2 .lut_mask = 64'h0660066006600660;
defparam \aneb_result_wire[0]~2 .shared_arith = "off";

endmodule

module Computer_System_dffpipe_3dc (
	dffe13a_0,
	clrn,
	clock)/* synthesis synthesis_greybox=0 */;
output 	dffe13a_0;
input 	clrn;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffe12a[0]~q ;


dffeas \dffe13a[0] (
	.clk(clock),
	.d(\dffe12a[0]~q ),
	.asdata(vcc),
	.clrn(!clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe13a_0),
	.prn(vcc));
defparam \dffe13a[0] .is_wysiwyg = "true";
defparam \dffe13a[0] .power_up = "low";

dffeas \dffe12a[0] (
	.clk(clock),
	.d(vcc),
	.asdata(vcc),
	.clrn(!clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe12a[0]~q ),
	.prn(vcc));
defparam \dffe12a[0] .is_wysiwyg = "true";
defparam \dffe12a[0] .power_up = "low";

endmodule

module Computer_System_dffpipe_3dc_1 (
	clock,
	dffe13a_0,
	clrn)/* synthesis synthesis_greybox=0 */;
input 	clock;
output 	dffe13a_0;
input 	clrn;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dffe12a[0]~q ;


dffeas \dffe13a[0] (
	.clk(clock),
	.d(\dffe12a[0]~q ),
	.asdata(vcc),
	.clrn(!clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe13a_0),
	.prn(vcc));
defparam \dffe13a[0] .is_wysiwyg = "true";
defparam \dffe13a[0] .power_up = "low";

dffeas \dffe12a[0] (
	.clk(clock),
	.d(vcc),
	.asdata(vcc),
	.clrn(!clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dffe12a[0]~q ),
	.prn(vcc));
defparam \dffe12a[0] .is_wysiwyg = "true";
defparam \dffe12a[0] .power_up = "low";

endmodule

module Computer_System_dffpipe_gd9 (
	clrn,
	dffe14a_0,
	dffe14a_1,
	dffe14a_2,
	dffe14a_3,
	dffe14a_4,
	dffe14a_5,
	dffe14a_6,
	dffe14a_7,
	xor7,
	xor3,
	xor0,
	xor1,
	xor2,
	xor6,
	xor4,
	xor5,
	clock)/* synthesis synthesis_greybox=0 */;
input 	clrn;
output 	dffe14a_0;
output 	dffe14a_1;
output 	dffe14a_2;
output 	dffe14a_3;
output 	dffe14a_4;
output 	dffe14a_5;
output 	dffe14a_6;
output 	dffe14a_7;
input 	xor7;
input 	xor3;
input 	xor0;
input 	xor1;
input 	xor2;
input 	xor6;
input 	xor4;
input 	xor5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \dffe14a[0] (
	.clk(clock),
	.d(xor0),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_0),
	.prn(vcc));
defparam \dffe14a[0] .is_wysiwyg = "true";
defparam \dffe14a[0] .power_up = "low";

dffeas \dffe14a[1] (
	.clk(clock),
	.d(xor1),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_1),
	.prn(vcc));
defparam \dffe14a[1] .is_wysiwyg = "true";
defparam \dffe14a[1] .power_up = "low";

dffeas \dffe14a[2] (
	.clk(clock),
	.d(xor2),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_2),
	.prn(vcc));
defparam \dffe14a[2] .is_wysiwyg = "true";
defparam \dffe14a[2] .power_up = "low";

dffeas \dffe14a[3] (
	.clk(clock),
	.d(xor3),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_3),
	.prn(vcc));
defparam \dffe14a[3] .is_wysiwyg = "true";
defparam \dffe14a[3] .power_up = "low";

dffeas \dffe14a[4] (
	.clk(clock),
	.d(xor4),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_4),
	.prn(vcc));
defparam \dffe14a[4] .is_wysiwyg = "true";
defparam \dffe14a[4] .power_up = "low";

dffeas \dffe14a[5] (
	.clk(clock),
	.d(xor5),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_5),
	.prn(vcc));
defparam \dffe14a[5] .is_wysiwyg = "true";
defparam \dffe14a[5] .power_up = "low";

dffeas \dffe14a[6] (
	.clk(clock),
	.d(xor6),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_6),
	.prn(vcc));
defparam \dffe14a[6] .is_wysiwyg = "true";
defparam \dffe14a[6] .power_up = "low";

dffeas \dffe14a[7] (
	.clk(clock),
	.d(xor7),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_7),
	.prn(vcc));
defparam \dffe14a[7] .is_wysiwyg = "true";
defparam \dffe14a[7] .power_up = "low";

endmodule

module Computer_System_dffpipe_gd9_1 (
	clrn,
	dffe14a_0,
	dffe14a_1,
	dffe14a_2,
	dffe14a_3,
	dffe14a_4,
	dffe14a_5,
	dffe14a_6,
	dffe14a_7,
	xor7,
	xor3,
	xor0,
	xor1,
	xor2,
	xor6,
	xor4,
	xor5,
	clock)/* synthesis synthesis_greybox=0 */;
input 	clrn;
output 	dffe14a_0;
output 	dffe14a_1;
output 	dffe14a_2;
output 	dffe14a_3;
output 	dffe14a_4;
output 	dffe14a_5;
output 	dffe14a_6;
output 	dffe14a_7;
input 	xor7;
input 	xor3;
input 	xor0;
input 	xor1;
input 	xor2;
input 	xor6;
input 	xor4;
input 	xor5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \dffe14a[0] (
	.clk(clock),
	.d(xor0),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_0),
	.prn(vcc));
defparam \dffe14a[0] .is_wysiwyg = "true";
defparam \dffe14a[0] .power_up = "low";

dffeas \dffe14a[1] (
	.clk(clock),
	.d(xor1),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_1),
	.prn(vcc));
defparam \dffe14a[1] .is_wysiwyg = "true";
defparam \dffe14a[1] .power_up = "low";

dffeas \dffe14a[2] (
	.clk(clock),
	.d(xor2),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_2),
	.prn(vcc));
defparam \dffe14a[2] .is_wysiwyg = "true";
defparam \dffe14a[2] .power_up = "low";

dffeas \dffe14a[3] (
	.clk(clock),
	.d(xor3),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_3),
	.prn(vcc));
defparam \dffe14a[3] .is_wysiwyg = "true";
defparam \dffe14a[3] .power_up = "low";

dffeas \dffe14a[4] (
	.clk(clock),
	.d(xor4),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_4),
	.prn(vcc));
defparam \dffe14a[4] .is_wysiwyg = "true";
defparam \dffe14a[4] .power_up = "low";

dffeas \dffe14a[5] (
	.clk(clock),
	.d(xor5),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_5),
	.prn(vcc));
defparam \dffe14a[5] .is_wysiwyg = "true";
defparam \dffe14a[5] .power_up = "low";

dffeas \dffe14a[6] (
	.clk(clock),
	.d(xor6),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_6),
	.prn(vcc));
defparam \dffe14a[6] .is_wysiwyg = "true";
defparam \dffe14a[6] .power_up = "low";

dffeas \dffe14a[7] (
	.clk(clock),
	.d(xor7),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_7),
	.prn(vcc));
defparam \dffe14a[7] .is_wysiwyg = "true";
defparam \dffe14a[7] .power_up = "low";

endmodule

module Computer_System_dffpipe_gd9_2 (
	clock,
	clrn,
	dffe14a_2,
	dffe14a_3,
	dffe14a_4,
	dffe14a_5,
	dffe14a_0,
	dffe14a_1,
	dffe14a_6,
	dffe14a_7,
	xor7,
	xor6,
	xor5,
	xor4,
	xor3,
	xor2,
	xor1,
	xor0)/* synthesis synthesis_greybox=0 */;
input 	clock;
input 	clrn;
output 	dffe14a_2;
output 	dffe14a_3;
output 	dffe14a_4;
output 	dffe14a_5;
output 	dffe14a_0;
output 	dffe14a_1;
output 	dffe14a_6;
output 	dffe14a_7;
input 	xor7;
input 	xor6;
input 	xor5;
input 	xor4;
input 	xor3;
input 	xor2;
input 	xor1;
input 	xor0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \dffe14a[2] (
	.clk(clock),
	.d(xor2),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_2),
	.prn(vcc));
defparam \dffe14a[2] .is_wysiwyg = "true";
defparam \dffe14a[2] .power_up = "low";

dffeas \dffe14a[3] (
	.clk(clock),
	.d(xor3),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_3),
	.prn(vcc));
defparam \dffe14a[3] .is_wysiwyg = "true";
defparam \dffe14a[3] .power_up = "low";

dffeas \dffe14a[4] (
	.clk(clock),
	.d(xor4),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_4),
	.prn(vcc));
defparam \dffe14a[4] .is_wysiwyg = "true";
defparam \dffe14a[4] .power_up = "low";

dffeas \dffe14a[5] (
	.clk(clock),
	.d(xor5),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_5),
	.prn(vcc));
defparam \dffe14a[5] .is_wysiwyg = "true";
defparam \dffe14a[5] .power_up = "low";

dffeas \dffe14a[0] (
	.clk(clock),
	.d(xor0),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_0),
	.prn(vcc));
defparam \dffe14a[0] .is_wysiwyg = "true";
defparam \dffe14a[0] .power_up = "low";

dffeas \dffe14a[1] (
	.clk(clock),
	.d(xor1),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_1),
	.prn(vcc));
defparam \dffe14a[1] .is_wysiwyg = "true";
defparam \dffe14a[1] .power_up = "low";

dffeas \dffe14a[6] (
	.clk(clock),
	.d(xor6),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_6),
	.prn(vcc));
defparam \dffe14a[6] .is_wysiwyg = "true";
defparam \dffe14a[6] .power_up = "low";

dffeas \dffe14a[7] (
	.clk(clock),
	.d(xor7),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_7),
	.prn(vcc));
defparam \dffe14a[7] .is_wysiwyg = "true";
defparam \dffe14a[7] .power_up = "low";

endmodule

module Computer_System_dffpipe_gd9_3 (
	clock,
	clrn,
	ram_address_a_7,
	dffe14a_2,
	dffe14a_3,
	dffe14a_4,
	dffe14a_5,
	dffe14a_0,
	dffe14a_1,
	dffe14a_6,
	dffe14a_7,
	xor6,
	xor5,
	xor4,
	xor3,
	xor2,
	xor1,
	xor0)/* synthesis synthesis_greybox=0 */;
input 	clock;
input 	clrn;
input 	ram_address_a_7;
output 	dffe14a_2;
output 	dffe14a_3;
output 	dffe14a_4;
output 	dffe14a_5;
output 	dffe14a_0;
output 	dffe14a_1;
output 	dffe14a_6;
output 	dffe14a_7;
input 	xor6;
input 	xor5;
input 	xor4;
input 	xor3;
input 	xor2;
input 	xor1;
input 	xor0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \dffe14a[2] (
	.clk(clock),
	.d(xor2),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_2),
	.prn(vcc));
defparam \dffe14a[2] .is_wysiwyg = "true";
defparam \dffe14a[2] .power_up = "low";

dffeas \dffe14a[3] (
	.clk(clock),
	.d(xor3),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_3),
	.prn(vcc));
defparam \dffe14a[3] .is_wysiwyg = "true";
defparam \dffe14a[3] .power_up = "low";

dffeas \dffe14a[4] (
	.clk(clock),
	.d(xor4),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_4),
	.prn(vcc));
defparam \dffe14a[4] .is_wysiwyg = "true";
defparam \dffe14a[4] .power_up = "low";

dffeas \dffe14a[5] (
	.clk(clock),
	.d(xor5),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_5),
	.prn(vcc));
defparam \dffe14a[5] .is_wysiwyg = "true";
defparam \dffe14a[5] .power_up = "low";

dffeas \dffe14a[0] (
	.clk(clock),
	.d(xor0),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_0),
	.prn(vcc));
defparam \dffe14a[0] .is_wysiwyg = "true";
defparam \dffe14a[0] .power_up = "low";

dffeas \dffe14a[1] (
	.clk(clock),
	.d(xor1),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_1),
	.prn(vcc));
defparam \dffe14a[1] .is_wysiwyg = "true";
defparam \dffe14a[1] .power_up = "low";

dffeas \dffe14a[6] (
	.clk(clock),
	.d(xor6),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_6),
	.prn(vcc));
defparam \dffe14a[6] .is_wysiwyg = "true";
defparam \dffe14a[6] .power_up = "low";

dffeas \dffe14a[7] (
	.clk(clock),
	.d(ram_address_a_7),
	.asdata(vcc),
	.clrn(clrn),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe14a_7),
	.prn(vcc));
defparam \dffe14a[7] .is_wysiwyg = "true";
defparam \dffe14a[7] .power_up = "low";

endmodule

module Computer_System_Computer_System_mm_interconnect_0 (
	h2f_ARVALID_0,
	h2f_AWVALID_0,
	h2f_BREADY_0,
	h2f_RREADY_0,
	h2f_WLAST_0,
	h2f_WVALID_0,
	h2f_ARADDR_0,
	h2f_ARADDR_1,
	h2f_ARADDR_2,
	h2f_ARADDR_3,
	h2f_ARADDR_4,
	h2f_ARADDR_5,
	h2f_ARADDR_6,
	h2f_ARADDR_7,
	h2f_ARADDR_8,
	h2f_ARADDR_9,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARLEN_0,
	h2f_ARLEN_1,
	h2f_ARLEN_2,
	h2f_ARLEN_3,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWADDR_0,
	h2f_AWADDR_1,
	h2f_AWADDR_2,
	h2f_AWADDR_3,
	h2f_AWADDR_4,
	h2f_AWADDR_5,
	h2f_AWADDR_6,
	h2f_AWADDR_7,
	h2f_AWADDR_8,
	h2f_AWADDR_9,
	h2f_AWADDR_10,
	h2f_AWADDR_11,
	h2f_AWADDR_12,
	h2f_AWADDR_13,
	h2f_AWADDR_14,
	h2f_AWADDR_15,
	h2f_AWADDR_16,
	h2f_AWADDR_17,
	h2f_AWADDR_18,
	h2f_AWADDR_19,
	h2f_AWADDR_20,
	h2f_AWADDR_21,
	h2f_AWADDR_22,
	h2f_AWADDR_23,
	h2f_AWADDR_24,
	h2f_AWADDR_25,
	h2f_AWADDR_26,
	h2f_AWADDR_27,
	h2f_AWBURST_0,
	h2f_AWBURST_1,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWLEN_0,
	h2f_AWLEN_1,
	h2f_AWLEN_2,
	h2f_AWLEN_3,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WDATA_1,
	h2f_WDATA_2,
	h2f_WDATA_3,
	h2f_WDATA_4,
	h2f_WDATA_5,
	h2f_WDATA_6,
	h2f_WDATA_7,
	h2f_WDATA_8,
	h2f_WDATA_9,
	h2f_WDATA_10,
	h2f_WDATA_11,
	h2f_WDATA_12,
	h2f_WDATA_13,
	h2f_WDATA_14,
	h2f_WDATA_15,
	h2f_WDATA_16,
	h2f_WDATA_17,
	h2f_WDATA_18,
	h2f_WDATA_19,
	h2f_WDATA_20,
	h2f_WDATA_21,
	h2f_WDATA_22,
	h2f_WDATA_23,
	h2f_WDATA_24,
	h2f_WDATA_25,
	h2f_WDATA_26,
	h2f_WDATA_27,
	h2f_WDATA_28,
	h2f_WDATA_29,
	h2f_WDATA_30,
	h2f_WDATA_31,
	h2f_WDATA_32,
	h2f_WDATA_33,
	h2f_WDATA_34,
	h2f_WDATA_35,
	h2f_WDATA_36,
	h2f_WDATA_37,
	h2f_WDATA_38,
	h2f_WDATA_39,
	h2f_WDATA_40,
	h2f_WDATA_41,
	h2f_WDATA_42,
	h2f_WDATA_43,
	h2f_WDATA_44,
	h2f_WDATA_45,
	h2f_WDATA_46,
	h2f_WDATA_47,
	h2f_WDATA_48,
	h2f_WDATA_49,
	h2f_WDATA_50,
	h2f_WDATA_51,
	h2f_WDATA_52,
	h2f_WDATA_53,
	h2f_WDATA_54,
	h2f_WDATA_55,
	h2f_WDATA_56,
	h2f_WDATA_57,
	h2f_WDATA_58,
	h2f_WDATA_59,
	h2f_WDATA_60,
	h2f_WDATA_61,
	h2f_WDATA_62,
	h2f_WDATA_63,
	h2f_WDATA_64,
	h2f_WDATA_65,
	h2f_WDATA_66,
	h2f_WDATA_67,
	h2f_WDATA_68,
	h2f_WDATA_69,
	h2f_WDATA_70,
	h2f_WDATA_71,
	h2f_WDATA_72,
	h2f_WDATA_73,
	h2f_WDATA_74,
	h2f_WDATA_75,
	h2f_WDATA_76,
	h2f_WDATA_77,
	h2f_WDATA_78,
	h2f_WDATA_79,
	h2f_WDATA_80,
	h2f_WDATA_81,
	h2f_WDATA_82,
	h2f_WDATA_83,
	h2f_WDATA_84,
	h2f_WDATA_85,
	h2f_WDATA_86,
	h2f_WDATA_87,
	h2f_WDATA_88,
	h2f_WDATA_89,
	h2f_WDATA_90,
	h2f_WDATA_91,
	h2f_WDATA_92,
	h2f_WDATA_93,
	h2f_WDATA_94,
	h2f_WDATA_95,
	h2f_WDATA_96,
	h2f_WDATA_97,
	h2f_WDATA_98,
	h2f_WDATA_99,
	h2f_WDATA_100,
	h2f_WDATA_101,
	h2f_WDATA_102,
	h2f_WDATA_103,
	h2f_WDATA_104,
	h2f_WDATA_105,
	h2f_WDATA_106,
	h2f_WDATA_107,
	h2f_WDATA_108,
	h2f_WDATA_109,
	h2f_WDATA_110,
	h2f_WDATA_111,
	h2f_WDATA_112,
	h2f_WDATA_113,
	h2f_WDATA_114,
	h2f_WDATA_115,
	h2f_WDATA_116,
	h2f_WDATA_117,
	h2f_WDATA_118,
	h2f_WDATA_119,
	h2f_WDATA_120,
	h2f_WDATA_121,
	h2f_WDATA_122,
	h2f_WDATA_123,
	h2f_WDATA_124,
	h2f_WDATA_125,
	h2f_WDATA_126,
	h2f_WDATA_127,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	h2f_WSTRB_4,
	h2f_WSTRB_5,
	h2f_WSTRB_6,
	h2f_WSTRB_7,
	h2f_WSTRB_8,
	h2f_WSTRB_9,
	h2f_WSTRB_10,
	h2f_WSTRB_11,
	h2f_WSTRB_12,
	h2f_WSTRB_13,
	h2f_WSTRB_14,
	h2f_WSTRB_15,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	outclk_wire_0,
	op_2,
	op_21,
	op_22,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_5,
	int_nxt_addr_reg_dly_6,
	int_nxt_addr_reg_dly_7,
	int_nxt_addr_reg_dly_8,
	int_nxt_addr_reg_dly_9,
	in_ready_hold,
	source0_data_34,
	source0_data_32,
	source0_data_33,
	source0_data_35,
	sink1_ready,
	wrfull,
	wrfull1,
	wrfull2,
	ARM_A9_HPS_h2f_axi_master_awready,
	WideOr1,
	src_payload_0,
	WideOr11,
	ARM_A9_HPS_h2f_axi_master_wready,
	src_data_209,
	src_data_210,
	src_data_211,
	src_data_212,
	src_data_213,
	src_data_214,
	src_data_215,
	src_data_216,
	src_data_217,
	src_data_218,
	src_data_219,
	src_data_220,
	src_data_0,
	src_payload,
	src_data_2,
	src_data_3,
	src_payload1,
	src_data_5,
	src_payload2,
	src_data_7,
	src_payload3,
	src_data_9,
	src_data_10,
	src_data_11,
	src_data_12,
	src_payload4,
	src_data_14,
	src_data_15,
	src_data_16,
	src_payload5,
	src_data_18,
	src_data_19,
	src_payload6,
	src_data_21,
	src_payload7,
	src_data_23,
	src_payload8,
	src_data_25,
	src_data_26,
	src_data_27,
	src_data_28,
	src_payload9,
	src_data_30,
	src_data_31,
	src_data_32,
	src_payload10,
	src_data_34,
	src_data_35,
	src_payload11,
	src_data_37,
	src_payload12,
	src_data_39,
	src_payload13,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_payload14,
	src_data_46,
	src_data_47,
	src_data_48,
	src_payload15,
	src_data_50,
	src_data_51,
	src_payload16,
	src_data_53,
	src_payload17,
	src_data_55,
	src_payload18,
	src_data_57,
	src_data_58,
	src_data_59,
	src_data_60,
	src_payload19,
	src_data_62,
	src_data_63,
	src_data_64,
	src_payload20,
	src_data_66,
	src_data_67,
	src_payload21,
	src_data_69,
	src_payload22,
	src_data_71,
	src_payload23,
	src_data_73,
	src_data_74,
	src_data_75,
	src_data_76,
	src_payload24,
	src_data_78,
	src_data_79,
	src_data_80,
	src_payload25,
	src_data_82,
	src_data_83,
	src_payload26,
	src_data_85,
	src_payload27,
	src_data_87,
	src_payload28,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_payload29,
	src_data_94,
	src_data_95,
	src_data_96,
	src_payload30,
	src_data_98,
	src_data_99,
	src_payload31,
	src_data_101,
	src_payload32,
	src_data_103,
	src_payload33,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	src_payload34,
	src_data_110,
	src_data_111,
	src_data_112,
	src_payload35,
	src_data_114,
	src_data_115,
	src_payload36,
	src_data_117,
	src_payload37,
	src_data_119,
	src_payload38,
	src_data_121,
	src_data_122,
	src_data_123,
	src_data_124,
	src_payload39,
	src_data_126,
	src_data_127,
	src_data_2091,
	src_data_2101,
	src_data_2111,
	src_data_2121,
	src_data_2131,
	src_data_2141,
	src_data_2151,
	src_data_2161,
	src_data_2171,
	src_data_2181,
	src_data_2191,
	src_data_2201,
	m0_write,
	in_data_reg_0,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	m0_write1,
	in_data_reg_01,
	in_data_reg_110,
	in_data_reg_210,
	in_data_reg_32,
	in_data_reg_41,
	in_data_reg_51,
	in_data_reg_61,
	in_data_reg_71,
	in_data_reg_81,
	in_data_reg_91,
	in_data_reg_101,
	in_data_reg_111,
	in_data_reg_121,
	in_data_reg_131,
	in_data_reg_141,
	in_data_reg_151,
	in_data_reg_161,
	in_data_reg_171,
	in_data_reg_181,
	in_data_reg_191,
	in_data_reg_201,
	in_data_reg_211,
	in_data_reg_221,
	in_data_reg_231,
	in_data_reg_241,
	in_data_reg_251,
	in_data_reg_261,
	in_data_reg_271,
	in_data_reg_281,
	in_data_reg_291,
	in_data_reg_301,
	in_data_reg_311,
	r_sync_rst,
	altera_reset_synchronizer_int_chain_out,
	wrfull3,
	wrfull4)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_AWVALID_0;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	h2f_WLAST_0;
input 	h2f_WVALID_0;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_3;
input 	h2f_ARADDR_4;
input 	h2f_ARADDR_5;
input 	h2f_ARADDR_6;
input 	h2f_ARADDR_7;
input 	h2f_ARADDR_8;
input 	h2f_ARADDR_9;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARLEN_0;
input 	h2f_ARLEN_1;
input 	h2f_ARLEN_2;
input 	h2f_ARLEN_3;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWADDR_0;
input 	h2f_AWADDR_1;
input 	h2f_AWADDR_2;
input 	h2f_AWADDR_3;
input 	h2f_AWADDR_4;
input 	h2f_AWADDR_5;
input 	h2f_AWADDR_6;
input 	h2f_AWADDR_7;
input 	h2f_AWADDR_8;
input 	h2f_AWADDR_9;
input 	h2f_AWADDR_10;
input 	h2f_AWADDR_11;
input 	h2f_AWADDR_12;
input 	h2f_AWADDR_13;
input 	h2f_AWADDR_14;
input 	h2f_AWADDR_15;
input 	h2f_AWADDR_16;
input 	h2f_AWADDR_17;
input 	h2f_AWADDR_18;
input 	h2f_AWADDR_19;
input 	h2f_AWADDR_20;
input 	h2f_AWADDR_21;
input 	h2f_AWADDR_22;
input 	h2f_AWADDR_23;
input 	h2f_AWADDR_24;
input 	h2f_AWADDR_25;
input 	h2f_AWADDR_26;
input 	h2f_AWADDR_27;
input 	h2f_AWBURST_0;
input 	h2f_AWBURST_1;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWLEN_0;
input 	h2f_AWLEN_1;
input 	h2f_AWLEN_2;
input 	h2f_AWLEN_3;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WDATA_1;
input 	h2f_WDATA_2;
input 	h2f_WDATA_3;
input 	h2f_WDATA_4;
input 	h2f_WDATA_5;
input 	h2f_WDATA_6;
input 	h2f_WDATA_7;
input 	h2f_WDATA_8;
input 	h2f_WDATA_9;
input 	h2f_WDATA_10;
input 	h2f_WDATA_11;
input 	h2f_WDATA_12;
input 	h2f_WDATA_13;
input 	h2f_WDATA_14;
input 	h2f_WDATA_15;
input 	h2f_WDATA_16;
input 	h2f_WDATA_17;
input 	h2f_WDATA_18;
input 	h2f_WDATA_19;
input 	h2f_WDATA_20;
input 	h2f_WDATA_21;
input 	h2f_WDATA_22;
input 	h2f_WDATA_23;
input 	h2f_WDATA_24;
input 	h2f_WDATA_25;
input 	h2f_WDATA_26;
input 	h2f_WDATA_27;
input 	h2f_WDATA_28;
input 	h2f_WDATA_29;
input 	h2f_WDATA_30;
input 	h2f_WDATA_31;
input 	h2f_WDATA_32;
input 	h2f_WDATA_33;
input 	h2f_WDATA_34;
input 	h2f_WDATA_35;
input 	h2f_WDATA_36;
input 	h2f_WDATA_37;
input 	h2f_WDATA_38;
input 	h2f_WDATA_39;
input 	h2f_WDATA_40;
input 	h2f_WDATA_41;
input 	h2f_WDATA_42;
input 	h2f_WDATA_43;
input 	h2f_WDATA_44;
input 	h2f_WDATA_45;
input 	h2f_WDATA_46;
input 	h2f_WDATA_47;
input 	h2f_WDATA_48;
input 	h2f_WDATA_49;
input 	h2f_WDATA_50;
input 	h2f_WDATA_51;
input 	h2f_WDATA_52;
input 	h2f_WDATA_53;
input 	h2f_WDATA_54;
input 	h2f_WDATA_55;
input 	h2f_WDATA_56;
input 	h2f_WDATA_57;
input 	h2f_WDATA_58;
input 	h2f_WDATA_59;
input 	h2f_WDATA_60;
input 	h2f_WDATA_61;
input 	h2f_WDATA_62;
input 	h2f_WDATA_63;
input 	h2f_WDATA_64;
input 	h2f_WDATA_65;
input 	h2f_WDATA_66;
input 	h2f_WDATA_67;
input 	h2f_WDATA_68;
input 	h2f_WDATA_69;
input 	h2f_WDATA_70;
input 	h2f_WDATA_71;
input 	h2f_WDATA_72;
input 	h2f_WDATA_73;
input 	h2f_WDATA_74;
input 	h2f_WDATA_75;
input 	h2f_WDATA_76;
input 	h2f_WDATA_77;
input 	h2f_WDATA_78;
input 	h2f_WDATA_79;
input 	h2f_WDATA_80;
input 	h2f_WDATA_81;
input 	h2f_WDATA_82;
input 	h2f_WDATA_83;
input 	h2f_WDATA_84;
input 	h2f_WDATA_85;
input 	h2f_WDATA_86;
input 	h2f_WDATA_87;
input 	h2f_WDATA_88;
input 	h2f_WDATA_89;
input 	h2f_WDATA_90;
input 	h2f_WDATA_91;
input 	h2f_WDATA_92;
input 	h2f_WDATA_93;
input 	h2f_WDATA_94;
input 	h2f_WDATA_95;
input 	h2f_WDATA_96;
input 	h2f_WDATA_97;
input 	h2f_WDATA_98;
input 	h2f_WDATA_99;
input 	h2f_WDATA_100;
input 	h2f_WDATA_101;
input 	h2f_WDATA_102;
input 	h2f_WDATA_103;
input 	h2f_WDATA_104;
input 	h2f_WDATA_105;
input 	h2f_WDATA_106;
input 	h2f_WDATA_107;
input 	h2f_WDATA_108;
input 	h2f_WDATA_109;
input 	h2f_WDATA_110;
input 	h2f_WDATA_111;
input 	h2f_WDATA_112;
input 	h2f_WDATA_113;
input 	h2f_WDATA_114;
input 	h2f_WDATA_115;
input 	h2f_WDATA_116;
input 	h2f_WDATA_117;
input 	h2f_WDATA_118;
input 	h2f_WDATA_119;
input 	h2f_WDATA_120;
input 	h2f_WDATA_121;
input 	h2f_WDATA_122;
input 	h2f_WDATA_123;
input 	h2f_WDATA_124;
input 	h2f_WDATA_125;
input 	h2f_WDATA_126;
input 	h2f_WDATA_127;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
input 	h2f_WSTRB_4;
input 	h2f_WSTRB_5;
input 	h2f_WSTRB_6;
input 	h2f_WSTRB_7;
input 	h2f_WSTRB_8;
input 	h2f_WSTRB_9;
input 	h2f_WSTRB_10;
input 	h2f_WSTRB_11;
input 	h2f_WSTRB_12;
input 	h2f_WSTRB_13;
input 	h2f_WSTRB_14;
input 	h2f_WSTRB_15;
input 	q_b_0;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	q_b_8;
input 	q_b_9;
input 	q_b_10;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_20;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_24;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_28;
input 	q_b_29;
input 	q_b_30;
input 	q_b_31;
input 	outclk_wire_0;
input 	op_2;
input 	op_21;
input 	op_22;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_5;
output 	int_nxt_addr_reg_dly_6;
output 	int_nxt_addr_reg_dly_7;
output 	int_nxt_addr_reg_dly_8;
output 	int_nxt_addr_reg_dly_9;
input 	in_ready_hold;
output 	source0_data_34;
output 	source0_data_32;
output 	source0_data_33;
output 	source0_data_35;
output 	sink1_ready;
input 	wrfull;
input 	wrfull1;
input 	wrfull2;
output 	ARM_A9_HPS_h2f_axi_master_awready;
output 	WideOr1;
output 	src_payload_0;
output 	WideOr11;
output 	ARM_A9_HPS_h2f_axi_master_wready;
output 	src_data_209;
output 	src_data_210;
output 	src_data_211;
output 	src_data_212;
output 	src_data_213;
output 	src_data_214;
output 	src_data_215;
output 	src_data_216;
output 	src_data_217;
output 	src_data_218;
output 	src_data_219;
output 	src_data_220;
output 	src_data_0;
output 	src_payload;
output 	src_data_2;
output 	src_data_3;
output 	src_payload1;
output 	src_data_5;
output 	src_payload2;
output 	src_data_7;
output 	src_payload3;
output 	src_data_9;
output 	src_data_10;
output 	src_data_11;
output 	src_data_12;
output 	src_payload4;
output 	src_data_14;
output 	src_data_15;
output 	src_data_16;
output 	src_payload5;
output 	src_data_18;
output 	src_data_19;
output 	src_payload6;
output 	src_data_21;
output 	src_payload7;
output 	src_data_23;
output 	src_payload8;
output 	src_data_25;
output 	src_data_26;
output 	src_data_27;
output 	src_data_28;
output 	src_payload9;
output 	src_data_30;
output 	src_data_31;
output 	src_data_32;
output 	src_payload10;
output 	src_data_34;
output 	src_data_35;
output 	src_payload11;
output 	src_data_37;
output 	src_payload12;
output 	src_data_39;
output 	src_payload13;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_payload14;
output 	src_data_46;
output 	src_data_47;
output 	src_data_48;
output 	src_payload15;
output 	src_data_50;
output 	src_data_51;
output 	src_payload16;
output 	src_data_53;
output 	src_payload17;
output 	src_data_55;
output 	src_payload18;
output 	src_data_57;
output 	src_data_58;
output 	src_data_59;
output 	src_data_60;
output 	src_payload19;
output 	src_data_62;
output 	src_data_63;
output 	src_data_64;
output 	src_payload20;
output 	src_data_66;
output 	src_data_67;
output 	src_payload21;
output 	src_data_69;
output 	src_payload22;
output 	src_data_71;
output 	src_payload23;
output 	src_data_73;
output 	src_data_74;
output 	src_data_75;
output 	src_data_76;
output 	src_payload24;
output 	src_data_78;
output 	src_data_79;
output 	src_data_80;
output 	src_payload25;
output 	src_data_82;
output 	src_data_83;
output 	src_payload26;
output 	src_data_85;
output 	src_payload27;
output 	src_data_87;
output 	src_payload28;
output 	src_data_89;
output 	src_data_90;
output 	src_data_91;
output 	src_data_92;
output 	src_payload29;
output 	src_data_94;
output 	src_data_95;
output 	src_data_96;
output 	src_payload30;
output 	src_data_98;
output 	src_data_99;
output 	src_payload31;
output 	src_data_101;
output 	src_payload32;
output 	src_data_103;
output 	src_payload33;
output 	src_data_105;
output 	src_data_106;
output 	src_data_107;
output 	src_data_108;
output 	src_payload34;
output 	src_data_110;
output 	src_data_111;
output 	src_data_112;
output 	src_payload35;
output 	src_data_114;
output 	src_data_115;
output 	src_payload36;
output 	src_data_117;
output 	src_payload37;
output 	src_data_119;
output 	src_payload38;
output 	src_data_121;
output 	src_data_122;
output 	src_data_123;
output 	src_data_124;
output 	src_payload39;
output 	src_data_126;
output 	src_data_127;
output 	src_data_2091;
output 	src_data_2101;
output 	src_data_2111;
output 	src_data_2121;
output 	src_data_2131;
output 	src_data_2141;
output 	src_data_2151;
output 	src_data_2161;
output 	src_data_2171;
output 	src_data_2181;
output 	src_data_2191;
output 	src_data_2201;
output 	m0_write;
output 	in_data_reg_0;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
output 	m0_write1;
output 	in_data_reg_01;
output 	in_data_reg_110;
output 	in_data_reg_210;
output 	in_data_reg_32;
output 	in_data_reg_41;
output 	in_data_reg_51;
output 	in_data_reg_61;
output 	in_data_reg_71;
output 	in_data_reg_81;
output 	in_data_reg_91;
output 	in_data_reg_101;
output 	in_data_reg_111;
output 	in_data_reg_121;
output 	in_data_reg_131;
output 	in_data_reg_141;
output 	in_data_reg_151;
output 	in_data_reg_161;
output 	in_data_reg_171;
output 	in_data_reg_181;
output 	in_data_reg_191;
output 	in_data_reg_201;
output 	in_data_reg_211;
output 	in_data_reg_221;
output 	in_data_reg_231;
output 	in_data_reg_241;
output 	in_data_reg_251;
output 	in_data_reg_261;
output 	in_data_reg_271;
output 	in_data_reg_281;
output 	in_data_reg_291;
output 	in_data_reg_301;
output 	in_data_reg_311;
input 	r_sync_rst;
input 	altera_reset_synchronizer_int_chain_out;
input 	wrfull3;
input 	wrfull4;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[24]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[25]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[23]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[13]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[21]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[22]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[19]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[20]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[15]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[16]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[17]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[18]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[26]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[27]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[12]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[14]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[10]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[11]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[9]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[8]~q ;
wire \fifo_hps_to_fpga_in_rsp_width_adapter|data_reg[0]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[0]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[1]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[2]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[3]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[4]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[5]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[6]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[7]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[8]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[9]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[10]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[11]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[12]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[13]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[14]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[15]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[16]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[17]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[18]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[19]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[20]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[21]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[22]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[23]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[24]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[25]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[26]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[27]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[28]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[29]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[30]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[31]~q ;
wire \fifo_hps_to_fpga_in_rsp_width_adapter|data_reg[32]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[32]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[33]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[34]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[35]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[36]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[37]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[38]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[39]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[40]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[41]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[42]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[43]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[44]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[45]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[46]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[47]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[48]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[49]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[50]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[51]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[52]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[53]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[54]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[55]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[56]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[57]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[58]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[59]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[60]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[61]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[62]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[63]~q ;
wire \fifo_hps_to_fpga_in_rsp_width_adapter|data_reg[64]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[64]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[65]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[66]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[67]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[68]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[69]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[70]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[71]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[72]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[73]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[74]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[75]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[76]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[77]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[78]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[79]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[80]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[81]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[82]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[83]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[84]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[85]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[86]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[87]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[88]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[89]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[90]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[91]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[92]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[93]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[94]~q ;
wire \onchip_sram_s2_rsp_width_adapter|data_reg[95]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|Add4~1_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add5~1_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add4~5_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add5~5_sumout ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[7]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[8]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|Add4~9_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add5~9_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add4~13_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add5~13_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add4~17_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add5~17_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add5~21_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add4~21_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add5~25_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add4~25_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add4~29_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add5~29_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add4~33_sumout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add5~33_sumout ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[2]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[3]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[1]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[1]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[0]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[0]~q ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|out_data[37]~3_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux4~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux5~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux6~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux7~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux8~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux9~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux10~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux11~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux12~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux13~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux14~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux15~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux16~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux17~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux18~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux19~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux20~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux21~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux22~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux23~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux24~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux25~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux26~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux27~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux28~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux29~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux30~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux31~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux32~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux33~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux34~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux35~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux4~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux5~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux6~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux7~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux8~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux9~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux10~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux11~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux12~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux13~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux14~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux15~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux16~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux17~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux18~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux19~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux20~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux21~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux22~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux23~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux24~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux25~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux26~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux27~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux28~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux29~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux30~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux31~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux32~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux33~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux34~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux35~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux3~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux2~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux1~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|Mux0~0_combout ;
wire \cmd_mux_001|src_data[185]~43_combout ;
wire \cmd_mux_001|saved_grant[1]~q ;
wire \cmd_mux_001|saved_grant[0]~q ;
wire \cmd_mux_001|src_data[198]~combout ;
wire \cmd_mux_001|src_data[199]~combout ;
wire \cmd_mux_001|src_data[200]~combout ;
wire \onchip_sram_s2_cmd_width_adapter|in_ready~0_combout ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|always12~0_combout ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~3_combout ;
wire \onchip_sram_s2_agent_rsp_fifo|mem_used[1]~q ;
wire \onchip_sram_s2_agent|cp_ready~combout ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_eop_reg~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|new_burst_reg~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_bytecount_reg_zero~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|ShiftLeft1~0_combout ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~5_combout ;
wire \onchip_sram_s2_agent|WideOr0~0_combout ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|sop_enable~q ;
wire \router|Equal0~6_combout ;
wire \router|Equal0~7_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[7]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[6]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[2]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[3]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[4]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[5]~q ;
wire \router|Equal0~14_combout ;
wire \cmd_demux|sink_ready~0_combout ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \fifo_hps_to_fpga_in_agent|WideOr0~0_combout ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem_used[1]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|load_next_out_cmd~combout ;
wire \router|Equal0~16_combout ;
wire \cmd_mux|saved_grant[0]~q ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|count[1]~q ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|count[0]~q ;
wire \cmd_demux|sink_ready~2_combout ;
wire \arm_a9_hps_h2f_axi_master_wr_limiter|last_channel[0]~q ;
wire \arm_a9_hps_h2f_axi_master_wr_limiter|has_pending_responses~q ;
wire \arm_a9_hps_h2f_axi_master_wr_limiter|cmd_sink_ready~0_combout ;
wire \cmd_mux|last_cycle~0_combout ;
wire \onchip_sram_s2_translator|read_latency_shift_reg[0]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem_used[0]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][125]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem_used[0]~q ;
wire \onchip_sram_s2_rsp_width_adapter|out_valid~0_combout ;
wire \onchip_sram_s2_agent|comb~0_combout ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][126]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][66]~q ;
wire \onchip_sram_s2_agent|uncompressor|burst_uncompress_busy~q ;
wire \onchip_sram_s2_agent|uncompressor|last_packet_beat~0_combout ;
wire \onchip_sram_s2_agent|uncompressor|last_packet_beat~1_combout ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][80]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][79]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][78]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][77]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][76]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][75]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][74]~q ;
wire \onchip_sram_s2_agent|uncompressor|last_packet_beat~4_combout ;
wire \rsp_mux_001|src_payload~0_combout ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][38]~q ;
wire \onchip_sram_s2_agent|uncompressor|source_addr[2]~0_combout ;
wire \onchip_sram_s2_agent|uncompressor|source_addr[2]~1_combout ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][122]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][123]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][91]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][124]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][90]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][39]~q ;
wire \onchip_sram_s2_agent|uncompressor|source_addr[3]~2_combout ;
wire \onchip_sram_s2_rsp_width_adapter|always10~9_combout ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][68]~q ;
wire \rsp_demux_001|src0_valid~0_combout ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][68]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][125]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem_used[0]~q ;
wire \fifo_hps_to_fpga_in_agent|comb~0_combout ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][122]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][123]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][124]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][90]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][91]~q ;
wire \fifo_hps_to_fpga_in_rsp_width_adapter|ShiftRight0~0_combout ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][38]~q ;
wire \fifo_hps_to_fpga_in_agent|uncompressor|source_addr[2]~0_combout ;
wire \fifo_hps_to_fpga_in_rsp_width_adapter|always10~0_combout ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][126]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][39]~q ;
wire \fifo_hps_to_fpga_in_agent|uncompressor|source_addr[3]~1_combout ;
wire \fifo_hps_to_fpga_in_rsp_width_adapter|always10~1_combout ;
wire \rsp_demux|src0_valid~0_combout ;
wire \rsp_demux|src1_valid~0_combout ;
wire \cmd_mux|last_cycle~1_combout ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][101]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][101]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][102]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][102]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][103]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][103]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][104]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][104]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][105]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][105]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][106]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][106]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][107]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][107]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][108]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][108]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][109]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][109]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][110]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][110]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][111]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][111]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][112]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][112]~q ;
wire \fifo_hps_to_fpga_in_agent_rdata_fifo|mem[0][31]~q ;
wire \fifo_hps_to_fpga_in_rsp_width_adapter|LessThan15~0_combout ;
wire \onchip_sram_s2_rsp_width_adapter|ShiftLeft0~0_combout ;
wire \onchip_sram_s2_agent_rdata_fifo|always4~0_combout ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][0]~q ;
wire \onchip_sram_s2_rsp_width_adapter|LessThan15~0_combout ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][1]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][2]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][3]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][4]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][5]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][6]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][7]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][8]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][9]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][10]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][11]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][12]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][13]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][14]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][15]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][16]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][17]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][18]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][19]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][20]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][21]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][22]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][23]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][24]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][25]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][26]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][27]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][28]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][29]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][30]~q ;
wire \onchip_sram_s2_agent_rdata_fifo|mem[0][31]~q ;
wire \onchip_sram_s2_rsp_width_adapter|ShiftLeft0~1_combout ;
wire \onchip_sram_s2_rsp_width_adapter|ShiftLeft0~2_combout ;
wire \onchip_sram_s2_agent_rdata_fifo|out_data[1]~0_combout ;
wire \onchip_sram_s2_agent_rdata_fifo|out_data[4]~1_combout ;
wire \onchip_sram_s2_agent_rdata_fifo|out_data[6]~2_combout ;
wire \onchip_sram_s2_agent_rdata_fifo|out_data[8]~3_combout ;
wire \onchip_sram_s2_agent_rdata_fifo|out_data[13]~4_combout ;
wire \onchip_sram_s2_agent_rdata_fifo|out_data[17]~5_combout ;
wire \onchip_sram_s2_agent_rdata_fifo|out_data[20]~6_combout ;
wire \onchip_sram_s2_agent_rdata_fifo|out_data[22]~7_combout ;
wire \onchip_sram_s2_agent_rdata_fifo|out_data[24]~8_combout ;
wire \onchip_sram_s2_agent_rdata_fifo|out_data[29]~9_combout ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ;
wire \router|Equal0~17_combout ;
wire \arm_a9_hps_h2f_axi_master_rd_limiter|cmd_src_valid[1]~0_combout ;
wire \arm_a9_hps_h2f_axi_master_wr_limiter|last_channel[1]~q ;
wire \cmd_demux|src1_valid~0_combout ;
wire \cmd_mux_001|WideOr1~combout ;
wire \cmd_mux_001|src_payload[0]~combout ;
wire \onchip_sram_s2_cmd_width_adapter|use_reg~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ;
wire \onchip_sram_s2_cmd_width_adapter|out_data[91]~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|out_data[90]~1_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|LessThan11~0_combout ;
wire \cmd_mux_001|src_payload~0_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add3~0_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|log2ceil~0_combout ;
wire \cmd_mux_001|src_data[190]~1_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[1]~q ;
wire \onchip_sram_s2_cmd_width_adapter|out_data[37]~3_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|LessThan10~0_combout ;
wire \cmd_mux_001|src_payload~1_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add3~1_combout ;
wire \cmd_mux_001|src_data[189]~4_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[0]~q ;
wire \cmd_mux_001|src_data[144]~combout ;
wire \onchip_sram_s2_cmd_width_adapter|out_data[36]~4_combout ;
wire \cmd_mux_001|src_data[130]~combout ;
wire \cmd_mux_001|src_data[134]~combout ;
wire \cmd_mux_001|src_data[138]~combout ;
wire \cmd_mux_001|src_data[142]~combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[2]~0_combout ;
wire \cmd_mux_001|src_data[146]~combout ;
wire \onchip_sram_s2_cmd_width_adapter|int_output_sel[0]~0_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[3]~1_combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux1~0_combout ;
wire \cmd_mux_001|src_data[128]~combout ;
wire \cmd_mux_001|src_data[132]~combout ;
wire \cmd_mux_001|src_data[136]~combout ;
wire \cmd_mux_001|src_data[140]~combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux3~0_combout ;
wire \cmd_mux_001|src_data[129]~combout ;
wire \cmd_mux_001|src_data[133]~combout ;
wire \cmd_mux_001|src_data[137]~combout ;
wire \cmd_mux_001|src_data[141]~combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux2~0_combout ;
wire \cmd_mux_001|src_data[131]~combout ;
wire \cmd_mux_001|src_data[135]~combout ;
wire \cmd_mux_001|src_data[139]~combout ;
wire \cmd_mux_001|src_data[143]~combout ;
wire \onchip_sram_s2_cmd_width_adapter|Mux0~0_combout ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ;
wire \onchip_sram_s2_agent|uncompressor|last_packet_beat~5_combout ;
wire \onchip_sram_s2_rsp_width_adapter|p1_ready~0_combout ;
wire \onchip_sram_s2_agent|cp_ready~0_combout ;
wire \onchip_sram_s2_cmd_width_adapter|out_endofpacket~2_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|burst_bytecount[4]~q ;
wire \cmd_mux_001|src_data[184]~combout ;
wire \arm_a9_hps_h2f_axi_master_agent|burst_bytecount[6]~q ;
wire \cmd_mux_001|src_payload~2_combout ;
wire \cmd_mux_001|src_payload~3_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|burst_bytecount[5]~q ;
wire \cmd_mux_001|src_payload~4_combout ;
wire \cmd_mux_001|src_payload~5_combout ;
wire \onchip_sram_s2_cmd_width_adapter|out_data[74]~5_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|burst_bytecount[7]~q ;
wire \arm_a9_hps_h2f_axi_master_agent|Add0~0_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add2~0_combout ;
wire \cmd_mux_001|src_data[187]~combout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add0~1_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add2~1_combout ;
wire \cmd_mux_001|src_data[186]~combout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add2~2_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|write_cp_data[188]~0_combout ;
wire \cmd_mux_001|src_payload~6_combout ;
wire \cmd_mux_001|src_data[188]~combout ;
wire \onchip_sram_s2_cmd_width_adapter|out_data[79]~6_combout ;
wire \onchip_sram_s2_cmd_width_adapter|out_data[76]~7_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|write_cp_data[187]~1_combout ;
wire \cmd_mux_001|src_payload~7_combout ;
wire \onchip_sram_s2_cmd_width_adapter|out_data[77]~11_combout ;
wire \onchip_sram_s2_cmd_width_adapter|out_data[78]~14_combout ;
wire \onchip_sram_s2_cmd_width_adapter|out_data[80]~15_combout ;
wire \onchip_sram_s2_cmd_width_adapter|out_data[75]~16_combout ;
wire \onchip_sram_s2_agent|cp_ready~1_combout ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \cmd_mux_001|src_valid~1_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[7]~20_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add1~3_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[9]~21_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[6]~22_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|LessThan16~0_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[8]~23_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|LessThan12~0_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|Selector26~0_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[4]~24_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|LessThan14~0_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[5]~25_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|LessThan15~0_combout ;
wire \cmd_demux|src0_valid~0_combout ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_eop_reg~q ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|LessThan2~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|int_output_sel[0]~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|int_output_sel[1]~1_combout ;
wire \fifo_hps_to_fpga_in_agent|cp_ready~0_combout ;
wire \fifo_hps_to_fpga_in_rsp_width_adapter|p1_ready~0_combout ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|read~0_combout ;
wire \cmd_mux|src_payload~0_combout ;
wire \cmd_mux|src_payload~1_combout ;
wire \cmd_mux|src_payload~2_combout ;
wire \fifo_hps_to_fpga_in_agent|cp_ready~1_combout ;
wire \cmd_demux|sink_ready~3_combout ;
wire \onchip_sram_s2_agent|WideOr0~combout ;
wire \onchip_sram_s2_rsp_width_adapter|always10~10_combout ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][83]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[122]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[123]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[124]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][84]~q ;
wire \fifo_hps_to_fpga_in_rsp_width_adapter|always10~2_combout ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[122]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[123]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[124]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][83]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][84]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[104]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[104]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ;
wire \cmd_mux_001|src_payload~8_combout ;
wire \cmd_mux_001|src_data[191]~6_combout ;
wire \cmd_mux_001|src_payload~9_combout ;
wire \cmd_mux_001|src_data[192]~7_combout ;
wire \cmd_mux_001|src_data[193]~8_combout ;
wire \cmd_mux_001|src_data[193]~10_combout ;
wire \onchip_sram_s2_cmd_width_adapter|address_reg[4]~q ;
wire \cmd_mux_001|src_payload~10_combout ;
wire \cmd_mux_001|src_data[194]~12_combout ;
wire \cmd_mux_001|src_data[194]~13_combout ;
wire \onchip_sram_s2_cmd_width_adapter|address_reg[5]~q ;
wire \cmd_mux_001|src_payload~11_combout ;
wire \cmd_mux_001|src_data[195]~15_combout ;
wire \cmd_mux_001|src_data[195]~16_combout ;
wire \onchip_sram_s2_cmd_width_adapter|address_reg[6]~q ;
wire \cmd_mux_001|src_payload~12_combout ;
wire \cmd_mux_001|src_data[196]~17_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|Add3~2_combout ;
wire \cmd_mux_001|src_data[196]~18_combout ;
wire \onchip_sram_s2_cmd_width_adapter|address_reg[7]~q ;
wire \cmd_mux_001|src_payload~13_combout ;
wire \cmd_mux_001|src_data[197]~19_combout ;
wire \cmd_mux_001|src_data[197]~20_combout ;
wire \cmd_mux_001|src_data[152]~combout ;
wire \onchip_sram_s2_cmd_width_adapter|out_data[44]~17_combout ;
wire \cmd_mux_001|src_payload~14_combout ;
wire \cmd_mux_001|src_payload~15_combout ;
wire \onchip_sram_s2_cmd_width_adapter|out_data[45]~18_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|Selector7~0_combout ;
wire \cmd_mux_001|src_data[190]~22_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[1]~26_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|Decoder0~1_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|Selector8~0_combout ;
wire \cmd_mux_001|src_data[189]~24_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[0]~27_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|out_endofpacket~1_combout ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ;
wire \cmd_demux|src0_valid~1_combout ;
wire \cmd_demux|sink_ready~4_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|out_data[90]~0_combout ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|out_data[91]~1_combout ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[2]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[3]~q ;
wire \cmd_mux|src_payload~3_combout ;
wire \cmd_mux_001|src_data[209]~combout ;
wire \cmd_mux|src_payload~4_combout ;
wire \cmd_mux_001|src_data[210]~combout ;
wire \cmd_mux|src_payload~5_combout ;
wire \cmd_mux_001|src_data[211]~combout ;
wire \cmd_mux|src_payload~6_combout ;
wire \cmd_mux_001|src_data[212]~combout ;
wire \cmd_mux|src_payload~7_combout ;
wire \cmd_mux_001|src_data[213]~combout ;
wire \cmd_mux|src_payload~8_combout ;
wire \cmd_mux_001|src_data[214]~combout ;
wire \cmd_mux|src_payload~9_combout ;
wire \cmd_mux_001|src_data[215]~combout ;
wire \cmd_mux|src_payload~10_combout ;
wire \cmd_mux_001|src_data[216]~combout ;
wire \cmd_mux|src_payload~11_combout ;
wire \cmd_mux_001|src_data[217]~combout ;
wire \cmd_mux|src_payload~12_combout ;
wire \cmd_mux_001|src_data[218]~combout ;
wire \cmd_mux|src_payload~13_combout ;
wire \cmd_mux_001|src_data[219]~combout ;
wire \cmd_mux|src_payload~14_combout ;
wire \cmd_mux_001|src_data[220]~combout ;
wire \arm_a9_hps_h2f_axi_master_agent|Selector6~0_combout ;
wire \cmd_mux_001|src_data[191]~26_combout ;
wire \arm_a9_hps_h2f_axi_master_agent|Selector5~0_combout ;
wire \cmd_mux_001|src_data[192]~28_combout ;
wire \cmd_mux_001|src_data[193]~31_combout ;
wire \cmd_mux_001|src_data[194]~34_combout ;
wire \cmd_mux_001|src_data[195]~37_combout ;
wire \cmd_mux_001|src_data[196]~40_combout ;
wire \cmd_mux_001|src_data[197]~42_combout ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][37]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][37]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][82]~q ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][36]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[1]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][82]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][36]~q ;
wire \fifo_hps_to_fpga_in_cmd_width_adapter|out_data[36]~2_combout ;
wire \onchip_sram_s2_agent_rsp_fifo|mem[0][81]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[1]~q ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[0]~q ;
wire \fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][81]~q ;
wire \cmd_mux|src_payload~15_combout ;
wire \fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[0]~q ;
wire \onchip_sram_s2_cmd_width_adapter|int_output_sel[1]~2_combout ;
wire \rsp_mux_001|src_payload~93_combout ;


Computer_System_Computer_System_mm_interconnect_0_cmd_mux_1 cmd_mux_001(
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_ARADDR_0(h2f_ARADDR_0),
	.h2f_ARADDR_2(h2f_ARADDR_2),
	.h2f_ARADDR_4(h2f_ARADDR_4),
	.h2f_ARADDR_5(h2f_ARADDR_5),
	.h2f_ARADDR_6(h2f_ARADDR_6),
	.h2f_ARADDR_7(h2f_ARADDR_7),
	.h2f_ARADDR_8(h2f_ARADDR_8),
	.h2f_ARADDR_9(h2f_ARADDR_9),
	.h2f_ARBURST_0(h2f_ARBURST_0),
	.h2f_ARBURST_1(h2f_ARBURST_1),
	.h2f_ARID_0(h2f_ARID_0),
	.h2f_ARID_1(h2f_ARID_1),
	.h2f_ARID_2(h2f_ARID_2),
	.h2f_ARID_3(h2f_ARID_3),
	.h2f_ARID_4(h2f_ARID_4),
	.h2f_ARID_5(h2f_ARID_5),
	.h2f_ARID_6(h2f_ARID_6),
	.h2f_ARID_7(h2f_ARID_7),
	.h2f_ARID_8(h2f_ARID_8),
	.h2f_ARID_9(h2f_ARID_9),
	.h2f_ARID_10(h2f_ARID_10),
	.h2f_ARID_11(h2f_ARID_11),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.h2f_ARLEN_1(h2f_ARLEN_1),
	.h2f_ARLEN_2(h2f_ARLEN_2),
	.h2f_ARLEN_3(h2f_ARLEN_3),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWADDR_0(h2f_AWADDR_0),
	.h2f_AWBURST_0(h2f_AWBURST_0),
	.h2f_AWBURST_1(h2f_AWBURST_1),
	.h2f_AWID_0(h2f_AWID_0),
	.h2f_AWID_1(h2f_AWID_1),
	.h2f_AWID_2(h2f_AWID_2),
	.h2f_AWID_3(h2f_AWID_3),
	.h2f_AWID_4(h2f_AWID_4),
	.h2f_AWID_5(h2f_AWID_5),
	.h2f_AWID_6(h2f_AWID_6),
	.h2f_AWID_7(h2f_AWID_7),
	.h2f_AWID_8(h2f_AWID_8),
	.h2f_AWID_9(h2f_AWID_9),
	.h2f_AWID_10(h2f_AWID_10),
	.h2f_AWID_11(h2f_AWID_11),
	.h2f_AWLEN_0(h2f_AWLEN_0),
	.h2f_AWLEN_1(h2f_AWLEN_1),
	.h2f_AWLEN_2(h2f_AWLEN_2),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.h2f_WSTRB_0(h2f_WSTRB_0),
	.h2f_WSTRB_1(h2f_WSTRB_1),
	.h2f_WSTRB_2(h2f_WSTRB_2),
	.h2f_WSTRB_3(h2f_WSTRB_3),
	.h2f_WSTRB_4(h2f_WSTRB_4),
	.h2f_WSTRB_5(h2f_WSTRB_5),
	.h2f_WSTRB_6(h2f_WSTRB_6),
	.h2f_WSTRB_7(h2f_WSTRB_7),
	.h2f_WSTRB_8(h2f_WSTRB_8),
	.h2f_WSTRB_9(h2f_WSTRB_9),
	.h2f_WSTRB_10(h2f_WSTRB_10),
	.h2f_WSTRB_11(h2f_WSTRB_11),
	.h2f_WSTRB_12(h2f_WSTRB_12),
	.h2f_WSTRB_13(h2f_WSTRB_13),
	.h2f_WSTRB_14(h2f_WSTRB_14),
	.h2f_WSTRB_15(h2f_WSTRB_15),
	.outclk_wire_0(outclk_wire_0),
	.Add4(\arm_a9_hps_h2f_axi_master_agent|Add4~1_sumout ),
	.Add5(\arm_a9_hps_h2f_axi_master_agent|Add5~1_sumout ),
	.Add41(\arm_a9_hps_h2f_axi_master_agent|Add4~5_sumout ),
	.Add51(\arm_a9_hps_h2f_axi_master_agent|Add5~5_sumout ),
	.Add42(\arm_a9_hps_h2f_axi_master_agent|Add4~9_sumout ),
	.Add52(\arm_a9_hps_h2f_axi_master_agent|Add5~9_sumout ),
	.Add43(\arm_a9_hps_h2f_axi_master_agent|Add4~13_sumout ),
	.Add53(\arm_a9_hps_h2f_axi_master_agent|Add5~13_sumout ),
	.Add44(\arm_a9_hps_h2f_axi_master_agent|Add4~17_sumout ),
	.Add54(\arm_a9_hps_h2f_axi_master_agent|Add5~17_sumout ),
	.Add55(\arm_a9_hps_h2f_axi_master_agent|Add5~21_sumout ),
	.Add45(\arm_a9_hps_h2f_axi_master_agent|Add4~21_sumout ),
	.Add56(\arm_a9_hps_h2f_axi_master_agent|Add5~25_sumout ),
	.Add46(\arm_a9_hps_h2f_axi_master_agent|Add4~25_sumout ),
	.Add47(\arm_a9_hps_h2f_axi_master_agent|Add4~29_sumout ),
	.Add57(\arm_a9_hps_h2f_axi_master_agent|Add5~29_sumout ),
	.Add48(\arm_a9_hps_h2f_axi_master_agent|Add4~33_sumout ),
	.Add58(\arm_a9_hps_h2f_axi_master_agent|Add5~33_sumout ),
	.src_data_185(\cmd_mux_001|src_data[185]~43_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.saved_grant_0(\cmd_mux_001|saved_grant[0]~q ),
	.src_data_198(\cmd_mux_001|src_data[198]~combout ),
	.src_data_199(\cmd_mux_001|src_data[199]~combout ),
	.src_data_200(\cmd_mux_001|src_data[200]~combout ),
	.in_ready(\onchip_sram_s2_cmd_width_adapter|in_ready~0_combout ),
	.nxt_in_ready(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready1(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.sink1_ready1(sink1_ready),
	.nxt_in_ready2(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ),
	.sop_enable(\arm_a9_hps_h2f_axi_master_agent|sop_enable~q ),
	.Equal0(\router|Equal0~6_combout ),
	.Equal01(\router|Equal0~7_combout ),
	.Equal02(\router|Equal0~14_combout ),
	.r_sync_rst(r_sync_rst),
	.Equal03(\router|Equal0~17_combout ),
	.cmd_src_valid_1(\arm_a9_hps_h2f_axi_master_rd_limiter|cmd_src_valid[1]~0_combout ),
	.src1_valid(\cmd_demux|src1_valid~0_combout ),
	.WideOr11(\cmd_mux_001|WideOr1~combout ),
	.src_payload_0(\cmd_mux_001|src_payload[0]~combout ),
	.LessThan11(\arm_a9_hps_h2f_axi_master_agent|LessThan11~0_combout ),
	.src_payload(\cmd_mux_001|src_payload~0_combout ),
	.Add3(\arm_a9_hps_h2f_axi_master_agent|Add3~0_combout ),
	.log2ceil(\arm_a9_hps_h2f_axi_master_agent|log2ceil~0_combout ),
	.src_data_190(\cmd_mux_001|src_data[190]~1_combout ),
	.LessThan10(\arm_a9_hps_h2f_axi_master_agent|LessThan10~0_combout ),
	.src_payload1(\cmd_mux_001|src_payload~1_combout ),
	.Add31(\arm_a9_hps_h2f_axi_master_agent|Add3~1_combout ),
	.src_data_189(\cmd_mux_001|src_data[189]~4_combout ),
	.address_burst_0(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[0]~q ),
	.src_data_144(\cmd_mux_001|src_data[144]~combout ),
	.src_data_130(\cmd_mux_001|src_data[130]~combout ),
	.src_data_134(\cmd_mux_001|src_data[134]~combout ),
	.src_data_138(\cmd_mux_001|src_data[138]~combout ),
	.src_data_142(\cmd_mux_001|src_data[142]~combout ),
	.out_data_2(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[2]~0_combout ),
	.src_data_146(\cmd_mux_001|src_data[146]~combout ),
	.src_data_128(\cmd_mux_001|src_data[128]~combout ),
	.src_data_132(\cmd_mux_001|src_data[132]~combout ),
	.src_data_136(\cmd_mux_001|src_data[136]~combout ),
	.src_data_140(\cmd_mux_001|src_data[140]~combout ),
	.src_data_129(\cmd_mux_001|src_data[129]~combout ),
	.src_data_133(\cmd_mux_001|src_data[133]~combout ),
	.src_data_137(\cmd_mux_001|src_data[137]~combout ),
	.src_data_141(\cmd_mux_001|src_data[141]~combout ),
	.src_data_131(\cmd_mux_001|src_data[131]~combout ),
	.src_data_135(\cmd_mux_001|src_data[135]~combout ),
	.src_data_139(\cmd_mux_001|src_data[139]~combout ),
	.src_data_143(\cmd_mux_001|src_data[143]~combout ),
	.burst_bytecount_4(\arm_a9_hps_h2f_axi_master_agent|burst_bytecount[4]~q ),
	.src_data_184(\cmd_mux_001|src_data[184]~combout ),
	.burst_bytecount_6(\arm_a9_hps_h2f_axi_master_agent|burst_bytecount[6]~q ),
	.src_payload2(\cmd_mux_001|src_payload~2_combout ),
	.src_payload3(\cmd_mux_001|src_payload~3_combout ),
	.burst_bytecount_5(\arm_a9_hps_h2f_axi_master_agent|burst_bytecount[5]~q ),
	.src_payload4(\cmd_mux_001|src_payload~4_combout ),
	.src_payload5(\cmd_mux_001|src_payload~5_combout ),
	.burst_bytecount_7(\arm_a9_hps_h2f_axi_master_agent|burst_bytecount[7]~q ),
	.Add0(\arm_a9_hps_h2f_axi_master_agent|Add0~0_combout ),
	.Add2(\arm_a9_hps_h2f_axi_master_agent|Add2~0_combout ),
	.src_data_187(\cmd_mux_001|src_data[187]~combout ),
	.Add01(\arm_a9_hps_h2f_axi_master_agent|Add0~1_combout ),
	.Add21(\arm_a9_hps_h2f_axi_master_agent|Add2~1_combout ),
	.src_data_186(\cmd_mux_001|src_data[186]~combout ),
	.Add22(\arm_a9_hps_h2f_axi_master_agent|Add2~2_combout ),
	.write_cp_data_188(\arm_a9_hps_h2f_axi_master_agent|write_cp_data[188]~0_combout ),
	.src_payload6(\cmd_mux_001|src_payload~6_combout ),
	.src_data_188(\cmd_mux_001|src_data[188]~combout ),
	.src_payload7(\cmd_mux_001|src_payload~7_combout ),
	.src_valid(\cmd_mux_001|src_valid~1_combout ),
	.Add1(\arm_a9_hps_h2f_axi_master_agent|Add1~3_combout ),
	.out_data_9(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[9]~21_combout ),
	.LessThan16(\arm_a9_hps_h2f_axi_master_agent|LessThan16~0_combout ),
	.out_data_8(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[8]~23_combout ),
	.LessThan12(\arm_a9_hps_h2f_axi_master_agent|LessThan12~0_combout ),
	.Selector26(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|Selector26~0_combout ),
	.LessThan14(\arm_a9_hps_h2f_axi_master_agent|LessThan14~0_combout ),
	.LessThan15(\arm_a9_hps_h2f_axi_master_agent|LessThan15~0_combout ),
	.src_payload8(\cmd_mux_001|src_payload~8_combout ),
	.src_data_191(\cmd_mux_001|src_data[191]~6_combout ),
	.src_payload9(\cmd_mux_001|src_payload~9_combout ),
	.src_data_192(\cmd_mux_001|src_data[192]~7_combout ),
	.src_data_193(\cmd_mux_001|src_data[193]~8_combout ),
	.src_data_1931(\cmd_mux_001|src_data[193]~10_combout ),
	.src_payload10(\cmd_mux_001|src_payload~10_combout ),
	.src_data_194(\cmd_mux_001|src_data[194]~12_combout ),
	.src_data_1941(\cmd_mux_001|src_data[194]~13_combout ),
	.src_payload11(\cmd_mux_001|src_payload~11_combout ),
	.src_data_195(\cmd_mux_001|src_data[195]~15_combout ),
	.src_data_1951(\cmd_mux_001|src_data[195]~16_combout ),
	.src_payload12(\cmd_mux_001|src_payload~12_combout ),
	.src_data_196(\cmd_mux_001|src_data[196]~17_combout ),
	.Add32(\arm_a9_hps_h2f_axi_master_agent|Add3~2_combout ),
	.src_data_1961(\cmd_mux_001|src_data[196]~18_combout ),
	.src_payload13(\cmd_mux_001|src_payload~13_combout ),
	.src_data_197(\cmd_mux_001|src_data[197]~19_combout ),
	.src_data_1971(\cmd_mux_001|src_data[197]~20_combout ),
	.src_data_152(\cmd_mux_001|src_data[152]~combout ),
	.src_payload14(\cmd_mux_001|src_payload~14_combout ),
	.src_payload15(\cmd_mux_001|src_payload~15_combout ),
	.Selector7(\arm_a9_hps_h2f_axi_master_agent|Selector7~0_combout ),
	.src_data_1901(\cmd_mux_001|src_data[190]~22_combout ),
	.Selector8(\arm_a9_hps_h2f_axi_master_agent|Selector8~0_combout ),
	.src_data_1891(\cmd_mux_001|src_data[189]~24_combout ),
	.src_data_209(\cmd_mux_001|src_data[209]~combout ),
	.src_data_210(\cmd_mux_001|src_data[210]~combout ),
	.src_data_211(\cmd_mux_001|src_data[211]~combout ),
	.src_data_212(\cmd_mux_001|src_data[212]~combout ),
	.src_data_213(\cmd_mux_001|src_data[213]~combout ),
	.src_data_214(\cmd_mux_001|src_data[214]~combout ),
	.src_data_215(\cmd_mux_001|src_data[215]~combout ),
	.src_data_216(\cmd_mux_001|src_data[216]~combout ),
	.src_data_217(\cmd_mux_001|src_data[217]~combout ),
	.src_data_218(\cmd_mux_001|src_data[218]~combout ),
	.src_data_219(\cmd_mux_001|src_data[219]~combout ),
	.src_data_220(\cmd_mux_001|src_data[220]~combout ),
	.Selector6(\arm_a9_hps_h2f_axi_master_agent|Selector6~0_combout ),
	.src_data_1911(\cmd_mux_001|src_data[191]~26_combout ),
	.Selector5(\arm_a9_hps_h2f_axi_master_agent|Selector5~0_combout ),
	.src_data_1921(\cmd_mux_001|src_data[192]~28_combout ),
	.src_data_1932(\cmd_mux_001|src_data[193]~31_combout ),
	.src_data_1942(\cmd_mux_001|src_data[194]~34_combout ),
	.src_data_1952(\cmd_mux_001|src_data[195]~37_combout ),
	.src_data_1962(\cmd_mux_001|src_data[196]~40_combout ),
	.src_data_1972(\cmd_mux_001|src_data[197]~42_combout ));

Computer_System_Computer_System_mm_interconnect_0_cmd_mux cmd_mux(
	.h2f_AWVALID_0(h2f_AWVALID_0),
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_WVALID_0(h2f_WVALID_0),
	.h2f_AWID_0(h2f_AWID_0),
	.h2f_AWID_1(h2f_AWID_1),
	.h2f_AWID_2(h2f_AWID_2),
	.h2f_AWID_3(h2f_AWID_3),
	.h2f_AWID_4(h2f_AWID_4),
	.h2f_AWID_5(h2f_AWID_5),
	.h2f_AWID_6(h2f_AWID_6),
	.h2f_AWID_7(h2f_AWID_7),
	.h2f_AWID_8(h2f_AWID_8),
	.h2f_AWID_9(h2f_AWID_9),
	.h2f_AWID_10(h2f_AWID_10),
	.h2f_AWID_11(h2f_AWID_11),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.outclk_wire_0(outclk_wire_0),
	.in_ready_hold(in_ready_hold),
	.Equal0(\router|Equal0~6_combout ),
	.Equal01(\router|Equal0~7_combout ),
	.Equal02(\router|Equal0~14_combout ),
	.nxt_in_ready(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.load_next_out_cmd(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|load_next_out_cmd~combout ),
	.Equal03(\router|Equal0~16_combout ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.sink_ready(\cmd_demux|sink_ready~2_combout ),
	.last_channel_0(\arm_a9_hps_h2f_axi_master_wr_limiter|last_channel[0]~q ),
	.has_pending_responses(\arm_a9_hps_h2f_axi_master_wr_limiter|has_pending_responses~q ),
	.last_cycle(\cmd_mux|last_cycle~0_combout ),
	.last_cycle1(\cmd_mux|last_cycle~1_combout ),
	.r_sync_rst(r_sync_rst),
	.src0_valid(\cmd_demux|src0_valid~0_combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.src_payload1(\cmd_mux|src_payload~1_combout ),
	.src_payload2(\cmd_mux|src_payload~2_combout ),
	.Selector7(\arm_a9_hps_h2f_axi_master_agent|Selector7~0_combout ),
	.nxt_in_ready1(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready2(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.src0_valid1(\cmd_demux|src0_valid~1_combout ),
	.sink_ready1(\cmd_demux|sink_ready~4_combout ),
	.src_payload3(\cmd_mux|src_payload~3_combout ),
	.src_payload4(\cmd_mux|src_payload~4_combout ),
	.src_payload5(\cmd_mux|src_payload~5_combout ),
	.src_payload6(\cmd_mux|src_payload~6_combout ),
	.src_payload7(\cmd_mux|src_payload~7_combout ),
	.src_payload8(\cmd_mux|src_payload~8_combout ),
	.src_payload9(\cmd_mux|src_payload~9_combout ),
	.src_payload10(\cmd_mux|src_payload~10_combout ),
	.src_payload11(\cmd_mux|src_payload~11_combout ),
	.src_payload12(\cmd_mux|src_payload~12_combout ),
	.src_payload13(\cmd_mux|src_payload~13_combout ),
	.src_payload14(\cmd_mux|src_payload~14_combout ),
	.src_payload15(\cmd_mux|src_payload~15_combout ));

Computer_System_Computer_System_mm_interconnect_0_cmd_demux cmd_demux(
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.in_ready_hold(in_ready_hold),
	.saved_grant_0(\cmd_mux_001|saved_grant[0]~q ),
	.in_ready(\onchip_sram_s2_cmd_width_adapter|in_ready~0_combout ),
	.nxt_in_ready(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready1(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.Equal0(\router|Equal0~6_combout ),
	.Equal01(\router|Equal0~7_combout ),
	.Equal02(\router|Equal0~14_combout ),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.nxt_in_ready2(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.load_next_out_cmd(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|load_next_out_cmd~combout ),
	.Equal03(\router|Equal0~16_combout ),
	.saved_grant_01(\cmd_mux|saved_grant[0]~q ),
	.count_1(\fifo_hps_to_fpga_in_cmd_width_adapter|count[1]~q ),
	.count_0(\fifo_hps_to_fpga_in_cmd_width_adapter|count[0]~q ),
	.sink_ready1(\cmd_demux|sink_ready~2_combout ),
	.last_channel_0(\arm_a9_hps_h2f_axi_master_wr_limiter|last_channel[0]~q ),
	.has_pending_responses(\arm_a9_hps_h2f_axi_master_wr_limiter|has_pending_responses~q ),
	.last_cycle(\cmd_mux|last_cycle~1_combout ),
	.last_channel_1(\arm_a9_hps_h2f_axi_master_wr_limiter|last_channel[1]~q ),
	.src1_valid(\cmd_demux|src1_valid~0_combout ),
	.src0_valid(\cmd_demux|src0_valid~0_combout ),
	.sink_ready2(\cmd_demux|sink_ready~3_combout ),
	.src0_valid1(\cmd_demux|src0_valid~1_combout ),
	.sink_ready3(\cmd_demux|sink_ready~4_combout ));

Computer_System_altera_merlin_burst_adapter_1 onchip_sram_s2_burst_adapter(
	.outclk_wire_0(outclk_wire_0),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_4(int_nxt_addr_reg_dly_4),
	.int_nxt_addr_reg_dly_5(int_nxt_addr_reg_dly_5),
	.int_nxt_addr_reg_dly_6(int_nxt_addr_reg_dly_6),
	.int_nxt_addr_reg_dly_7(int_nxt_addr_reg_dly_7),
	.int_nxt_addr_reg_dly_8(int_nxt_addr_reg_dly_8),
	.int_nxt_addr_reg_dly_9(int_nxt_addr_reg_dly_9),
	.out_uncomp_byte_cnt_reg_6(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_2(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_3(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_7(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[7]~q ),
	.out_uncomp_byte_cnt_reg_4(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_8(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[8]~q ),
	.out_uncomp_byte_cnt_reg_5(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_burstwrap_reg_2(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[2]~q ),
	.out_burstwrap_reg_3(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[3]~q ),
	.out_addr_reg_1(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[1]~q ),
	.out_burstwrap_reg_1(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[1]~q ),
	.out_addr_reg_0(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[0]~q ),
	.out_burstwrap_reg_0(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[0]~q ),
	.Mux4(\onchip_sram_s2_cmd_width_adapter|Mux4~0_combout ),
	.Mux5(\onchip_sram_s2_cmd_width_adapter|Mux5~0_combout ),
	.Mux6(\onchip_sram_s2_cmd_width_adapter|Mux6~0_combout ),
	.Mux7(\onchip_sram_s2_cmd_width_adapter|Mux7~0_combout ),
	.Mux8(\onchip_sram_s2_cmd_width_adapter|Mux8~0_combout ),
	.Mux9(\onchip_sram_s2_cmd_width_adapter|Mux9~0_combout ),
	.Mux10(\onchip_sram_s2_cmd_width_adapter|Mux10~0_combout ),
	.Mux11(\onchip_sram_s2_cmd_width_adapter|Mux11~0_combout ),
	.Mux12(\onchip_sram_s2_cmd_width_adapter|Mux12~0_combout ),
	.Mux13(\onchip_sram_s2_cmd_width_adapter|Mux13~0_combout ),
	.Mux14(\onchip_sram_s2_cmd_width_adapter|Mux14~0_combout ),
	.Mux15(\onchip_sram_s2_cmd_width_adapter|Mux15~0_combout ),
	.Mux16(\onchip_sram_s2_cmd_width_adapter|Mux16~0_combout ),
	.Mux17(\onchip_sram_s2_cmd_width_adapter|Mux17~0_combout ),
	.Mux18(\onchip_sram_s2_cmd_width_adapter|Mux18~0_combout ),
	.Mux19(\onchip_sram_s2_cmd_width_adapter|Mux19~0_combout ),
	.Mux20(\onchip_sram_s2_cmd_width_adapter|Mux20~0_combout ),
	.Mux21(\onchip_sram_s2_cmd_width_adapter|Mux21~0_combout ),
	.Mux22(\onchip_sram_s2_cmd_width_adapter|Mux22~0_combout ),
	.Mux23(\onchip_sram_s2_cmd_width_adapter|Mux23~0_combout ),
	.Mux24(\onchip_sram_s2_cmd_width_adapter|Mux24~0_combout ),
	.Mux25(\onchip_sram_s2_cmd_width_adapter|Mux25~0_combout ),
	.Mux26(\onchip_sram_s2_cmd_width_adapter|Mux26~0_combout ),
	.Mux27(\onchip_sram_s2_cmd_width_adapter|Mux27~0_combout ),
	.Mux28(\onchip_sram_s2_cmd_width_adapter|Mux28~0_combout ),
	.Mux29(\onchip_sram_s2_cmd_width_adapter|Mux29~0_combout ),
	.Mux30(\onchip_sram_s2_cmd_width_adapter|Mux30~0_combout ),
	.Mux31(\onchip_sram_s2_cmd_width_adapter|Mux31~0_combout ),
	.Mux32(\onchip_sram_s2_cmd_width_adapter|Mux32~0_combout ),
	.Mux33(\onchip_sram_s2_cmd_width_adapter|Mux33~0_combout ),
	.Mux34(\onchip_sram_s2_cmd_width_adapter|Mux34~0_combout ),
	.Mux35(\onchip_sram_s2_cmd_width_adapter|Mux35~0_combout ),
	.in_ready_hold(in_ready_hold),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.saved_grant_0(\cmd_mux_001|saved_grant[0]~q ),
	.src_data_198(\cmd_mux_001|src_data[198]~combout ),
	.src_data_199(\cmd_mux_001|src_data[199]~combout ),
	.src_data_200(\cmd_mux_001|src_data[200]~combout ),
	.stateST_COMP_TRANS(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.in_narrow_reg(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.always12(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|always12~0_combout ),
	.in_data_reg_91(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.in_data_reg_90(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ),
	.in_byteen_reg_2(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.source0_data_34(source0_data_34),
	.in_byteen_reg_0(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.source0_data_32(source0_data_32),
	.in_byteen_reg_1(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.source0_data_33(source0_data_33),
	.in_byteen_reg_3(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.source0_data_35(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~3_combout ),
	.source0_data_351(source0_data_35),
	.mem_used_1(\onchip_sram_s2_agent_rsp_fifo|mem_used[1]~q ),
	.cp_ready(\onchip_sram_s2_agent|cp_ready~combout ),
	.in_eop_reg(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_eop_reg~q ),
	.new_burst_reg(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|new_burst_reg~q ),
	.in_bytecount_reg_zero(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_bytecount_reg_zero~q ),
	.nxt_in_ready(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.out_valid_reg(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.ShiftLeft1(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|ShiftLeft1~0_combout ),
	.source0_data_352(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~5_combout ),
	.WideOr0(\onchip_sram_s2_agent|WideOr0~0_combout ),
	.nxt_in_ready2(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ),
	.in_data_reg_68(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.in_data_reg_0(in_data_reg_01),
	.in_data_reg_1(in_data_reg_110),
	.in_data_reg_2(in_data_reg_210),
	.in_data_reg_3(in_data_reg_32),
	.in_data_reg_4(in_data_reg_41),
	.in_data_reg_5(in_data_reg_51),
	.in_data_reg_6(in_data_reg_61),
	.in_data_reg_7(in_data_reg_71),
	.in_data_reg_8(in_data_reg_81),
	.in_data_reg_9(in_data_reg_91),
	.in_data_reg_10(in_data_reg_101),
	.in_data_reg_11(in_data_reg_111),
	.in_data_reg_12(in_data_reg_121),
	.in_data_reg_13(in_data_reg_131),
	.in_data_reg_14(in_data_reg_141),
	.in_data_reg_15(in_data_reg_151),
	.in_data_reg_16(in_data_reg_161),
	.in_data_reg_17(in_data_reg_171),
	.in_data_reg_18(in_data_reg_181),
	.in_data_reg_19(in_data_reg_191),
	.in_data_reg_20(in_data_reg_201),
	.in_data_reg_21(in_data_reg_211),
	.in_data_reg_22(in_data_reg_221),
	.in_data_reg_23(in_data_reg_231),
	.in_data_reg_24(in_data_reg_241),
	.in_data_reg_25(in_data_reg_251),
	.in_data_reg_26(in_data_reg_261),
	.in_data_reg_27(in_data_reg_271),
	.in_data_reg_28(in_data_reg_281),
	.in_data_reg_29(in_data_reg_291),
	.in_data_reg_30(in_data_reg_301),
	.in_data_reg_31(in_data_reg_311),
	.r_sync_rst(r_sync_rst),
	.WideOr1(\cmd_mux_001|WideOr1~combout ),
	.use_reg(\onchip_sram_s2_cmd_width_adapter|use_reg~q ),
	.nxt_out_eop(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.out_data_91(\onchip_sram_s2_cmd_width_adapter|out_data[91]~0_combout ),
	.out_data_90(\onchip_sram_s2_cmd_width_adapter|out_data[90]~1_combout ),
	.src_payload(\cmd_mux_001|src_payload~0_combout ),
	.src_data_190(\cmd_mux_001|src_data[190]~1_combout ),
	.out_data_37(\onchip_sram_s2_cmd_width_adapter|out_data[37]~3_combout ),
	.src_payload1(\cmd_mux_001|src_payload~1_combout ),
	.src_data_189(\cmd_mux_001|src_data[189]~4_combout ),
	.out_data_36(\onchip_sram_s2_cmd_width_adapter|out_data[36]~4_combout ),
	.int_output_sel_0(\onchip_sram_s2_cmd_width_adapter|int_output_sel[0]~0_combout ),
	.Mux1(\onchip_sram_s2_cmd_width_adapter|Mux1~0_combout ),
	.Mux3(\onchip_sram_s2_cmd_width_adapter|Mux3~0_combout ),
	.Mux2(\onchip_sram_s2_cmd_width_adapter|Mux2~0_combout ),
	.Mux0(\onchip_sram_s2_cmd_width_adapter|Mux0~0_combout ),
	.in_data_reg_69(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.cp_ready1(\onchip_sram_s2_agent|cp_ready~0_combout ),
	.out_endofpacket(\onchip_sram_s2_cmd_width_adapter|out_endofpacket~2_combout ),
	.out_data_74(\onchip_sram_s2_cmd_width_adapter|out_data[74]~5_combout ),
	.out_data_79(\onchip_sram_s2_cmd_width_adapter|out_data[79]~6_combout ),
	.out_data_76(\onchip_sram_s2_cmd_width_adapter|out_data[76]~7_combout ),
	.out_data_77(\onchip_sram_s2_cmd_width_adapter|out_data[77]~11_combout ),
	.out_data_78(\onchip_sram_s2_cmd_width_adapter|out_data[78]~14_combout ),
	.out_data_80(\onchip_sram_s2_cmd_width_adapter|out_data[80]~15_combout ),
	.out_data_75(\onchip_sram_s2_cmd_width_adapter|out_data[75]~16_combout ),
	.cp_ready2(\onchip_sram_s2_agent|cp_ready~1_combout ),
	.out_byte_cnt_reg_2(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.src_valid(\cmd_mux_001|src_valid~1_combout ),
	.out_data_7(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[7]~20_combout ),
	.out_data_6(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[6]~22_combout ),
	.out_data_4(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[4]~24_combout ),
	.out_data_5(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[5]~25_combout ),
	.in_data_reg_122(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[122]~q ),
	.in_data_reg_123(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[123]~q ),
	.in_data_reg_124(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[124]~q ),
	.in_data_reg_101(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.in_data_reg_104(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[104]~q ),
	.in_data_reg_105(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.src_payload2(\cmd_mux_001|src_payload~8_combout ),
	.src_data_191(\cmd_mux_001|src_data[191]~6_combout ),
	.src_payload3(\cmd_mux_001|src_payload~9_combout ),
	.src_data_192(\cmd_mux_001|src_data[192]~7_combout ),
	.src_data_193(\cmd_mux_001|src_data[193]~8_combout ),
	.src_data_1931(\cmd_mux_001|src_data[193]~10_combout ),
	.address_reg_4(\onchip_sram_s2_cmd_width_adapter|address_reg[4]~q ),
	.src_payload4(\cmd_mux_001|src_payload~10_combout ),
	.src_data_194(\cmd_mux_001|src_data[194]~12_combout ),
	.src_data_1941(\cmd_mux_001|src_data[194]~13_combout ),
	.address_reg_5(\onchip_sram_s2_cmd_width_adapter|address_reg[5]~q ),
	.src_payload5(\cmd_mux_001|src_payload~11_combout ),
	.src_data_195(\cmd_mux_001|src_data[195]~15_combout ),
	.src_data_1951(\cmd_mux_001|src_data[195]~16_combout ),
	.address_reg_6(\onchip_sram_s2_cmd_width_adapter|address_reg[6]~q ),
	.src_payload6(\cmd_mux_001|src_payload~12_combout ),
	.src_data_196(\cmd_mux_001|src_data[196]~17_combout ),
	.src_data_1961(\cmd_mux_001|src_data[196]~18_combout ),
	.address_reg_7(\onchip_sram_s2_cmd_width_adapter|address_reg[7]~q ),
	.src_payload7(\cmd_mux_001|src_payload~13_combout ),
	.src_data_197(\cmd_mux_001|src_data[197]~19_combout ),
	.src_data_1971(\cmd_mux_001|src_data[197]~20_combout ),
	.out_data_44(\onchip_sram_s2_cmd_width_adapter|out_data[44]~17_combout ),
	.out_data_45(\onchip_sram_s2_cmd_width_adapter|out_data[45]~18_combout ),
	.src_data_1901(\cmd_mux_001|src_data[190]~22_combout ),
	.src_data_1891(\cmd_mux_001|src_data[189]~24_combout ),
	.src_data_209(\cmd_mux_001|src_data[209]~combout ),
	.src_data_210(\cmd_mux_001|src_data[210]~combout ),
	.src_data_211(\cmd_mux_001|src_data[211]~combout ),
	.src_data_212(\cmd_mux_001|src_data[212]~combout ),
	.src_data_213(\cmd_mux_001|src_data[213]~combout ),
	.src_data_214(\cmd_mux_001|src_data[214]~combout ),
	.src_data_215(\cmd_mux_001|src_data[215]~combout ),
	.src_data_216(\cmd_mux_001|src_data[216]~combout ),
	.src_data_217(\cmd_mux_001|src_data[217]~combout ),
	.src_data_218(\cmd_mux_001|src_data[218]~combout ),
	.src_data_219(\cmd_mux_001|src_data[219]~combout ),
	.src_data_220(\cmd_mux_001|src_data[220]~combout ),
	.src_data_1911(\cmd_mux_001|src_data[191]~26_combout ),
	.src_data_1921(\cmd_mux_001|src_data[192]~28_combout ),
	.src_data_1932(\cmd_mux_001|src_data[193]~31_combout ),
	.src_data_1942(\cmd_mux_001|src_data[194]~34_combout ),
	.src_data_1952(\cmd_mux_001|src_data[195]~37_combout ),
	.src_data_1962(\cmd_mux_001|src_data[196]~40_combout ),
	.src_data_1972(\cmd_mux_001|src_data[197]~42_combout ),
	.int_output_sel_1(\onchip_sram_s2_cmd_width_adapter|int_output_sel[1]~2_combout ));

Computer_System_altera_merlin_burst_adapter fifo_hps_to_fpga_in_burst_adapter(
	.h2f_AWBURST_0(h2f_AWBURST_0),
	.h2f_AWBURST_1(h2f_AWBURST_1),
	.outclk_wire_0(outclk_wire_0),
	.Add4(\arm_a9_hps_h2f_axi_master_agent|Add4~9_sumout ),
	.Add41(\arm_a9_hps_h2f_axi_master_agent|Add4~13_sumout ),
	.out_data_37(\fifo_hps_to_fpga_in_cmd_width_adapter|out_data[37]~3_combout ),
	.Mux4(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux4~0_combout ),
	.Mux5(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux5~0_combout ),
	.Mux6(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux6~0_combout ),
	.Mux7(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux7~0_combout ),
	.Mux8(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux8~0_combout ),
	.Mux9(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux9~0_combout ),
	.Mux10(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux10~0_combout ),
	.Mux11(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux11~0_combout ),
	.Mux12(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux12~0_combout ),
	.Mux13(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux13~0_combout ),
	.Mux14(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux14~0_combout ),
	.Mux15(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux15~0_combout ),
	.Mux16(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux16~0_combout ),
	.Mux17(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux17~0_combout ),
	.Mux18(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux18~0_combout ),
	.Mux19(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux19~0_combout ),
	.Mux20(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux20~0_combout ),
	.Mux21(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux21~0_combout ),
	.Mux22(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux22~0_combout ),
	.Mux23(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux23~0_combout ),
	.Mux24(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux24~0_combout ),
	.Mux25(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux25~0_combout ),
	.Mux26(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux26~0_combout ),
	.Mux27(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux27~0_combout ),
	.Mux28(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux28~0_combout ),
	.Mux29(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux29~0_combout ),
	.Mux30(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux30~0_combout ),
	.Mux31(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux31~0_combout ),
	.Mux32(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux32~0_combout ),
	.Mux33(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux33~0_combout ),
	.Mux34(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux34~0_combout ),
	.Mux35(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux35~0_combout ),
	.Mux3(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux3~0_combout ),
	.Mux2(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux2~0_combout ),
	.Mux1(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux1~0_combout ),
	.Mux0(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux0~0_combout ),
	.in_ready_hold(in_ready_hold),
	.Equal0(\router|Equal0~6_combout ),
	.Equal01(\router|Equal0~7_combout ),
	.Equal02(\router|Equal0~14_combout ),
	.nxt_in_ready(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.out_valid_reg(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_byteen_reg_3(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\fifo_hps_to_fpga_in_agent|WideOr0~0_combout ),
	.wrfull(wrfull),
	.wrfull1(wrfull1),
	.wrfull2(wrfull2),
	.mem_used_1(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem_used[1]~q ),
	.load_next_out_cmd(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|load_next_out_cmd~combout ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.in_data_reg_68(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.nxt_uncomp_subburst_byte_cnt(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_uncomp_subburst_byte_cnt~0_combout ),
	.in_data_reg_0(in_data_reg_0),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_24(in_data_reg_24),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_31(in_data_reg_31),
	.r_sync_rst(r_sync_rst),
	.LessThan12(\arm_a9_hps_h2f_axi_master_agent|LessThan12~0_combout ),
	.Selector26(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|Selector26~0_combout ),
	.src0_valid(\cmd_demux|src0_valid~0_combout ),
	.in_eop_reg(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_eop_reg~q ),
	.wrfull3(wrfull3),
	.int_output_sel_0(\fifo_hps_to_fpga_in_cmd_width_adapter|int_output_sel[0]~0_combout ),
	.int_output_sel_1(\fifo_hps_to_fpga_in_cmd_width_adapter|int_output_sel[1]~1_combout ),
	.cp_ready(\fifo_hps_to_fpga_in_agent|cp_ready~0_combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.src_payload1(\cmd_mux|src_payload~1_combout ),
	.src_payload2(\cmd_mux|src_payload~2_combout ),
	.in_data_reg_122(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[122]~q ),
	.in_data_reg_123(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[123]~q ),
	.in_data_reg_124(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[124]~q ),
	.in_data_reg_90(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ),
	.in_data_reg_91(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.int_nxt_addr_reg_dly_2(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_3(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.in_data_reg_101(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.in_data_reg_104(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[104]~q ),
	.in_data_reg_105(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.Selector7(\arm_a9_hps_h2f_axi_master_agent|Selector7~0_combout ),
	.Selector8(\arm_a9_hps_h2f_axi_master_agent|Selector8~0_combout ),
	.out_endofpacket(\fifo_hps_to_fpga_in_cmd_width_adapter|out_endofpacket~1_combout ),
	.nxt_in_ready1(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready2(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.out_data_90(\fifo_hps_to_fpga_in_cmd_width_adapter|out_data[90]~0_combout ),
	.out_data_91(\fifo_hps_to_fpga_in_cmd_width_adapter|out_data[91]~1_combout ),
	.out_burstwrap_reg_2(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[2]~q ),
	.out_burstwrap_reg_3(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[3]~q ),
	.src_payload3(\cmd_mux|src_payload~3_combout ),
	.src_payload4(\cmd_mux|src_payload~4_combout ),
	.src_payload5(\cmd_mux|src_payload~5_combout ),
	.src_payload6(\cmd_mux|src_payload~6_combout ),
	.src_payload7(\cmd_mux|src_payload~7_combout ),
	.src_payload8(\cmd_mux|src_payload~8_combout ),
	.src_payload9(\cmd_mux|src_payload~9_combout ),
	.src_payload10(\cmd_mux|src_payload~10_combout ),
	.src_payload11(\cmd_mux|src_payload~11_combout ),
	.src_payload12(\cmd_mux|src_payload~12_combout ),
	.src_payload13(\cmd_mux|src_payload~13_combout ),
	.src_payload14(\cmd_mux|src_payload~14_combout ),
	.out_addr_reg_1(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[1]~q ),
	.out_data_36(\fifo_hps_to_fpga_in_cmd_width_adapter|out_data[36]~2_combout ),
	.out_burstwrap_reg_1(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[1]~q ),
	.out_addr_reg_0(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[0]~q ),
	.src_payload15(\cmd_mux|src_payload~15_combout ),
	.out_burstwrap_reg_0(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[0]~q ));

Computer_System_altera_merlin_traffic_limiter arm_a9_hps_h2f_axi_master_rd_limiter(
	.h2f_ARVALID_0(h2f_ARVALID_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.clk(outclk_wire_0),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.in_ready(\onchip_sram_s2_cmd_width_adapter|in_ready~0_combout ),
	.sink1_ready(sink1_ready),
	.nxt_in_ready(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ),
	.out_valid(\onchip_sram_s2_rsp_width_adapter|out_valid~0_combout ),
	.src_payload(\rsp_mux_001|src_payload~0_combout ),
	.src0_valid(\rsp_demux_001|src0_valid~0_combout ),
	.src_payload_0(src_payload_0),
	.WideOr1(WideOr11),
	.cmd_src_valid_1(\arm_a9_hps_h2f_axi_master_rd_limiter|cmd_src_valid[1]~0_combout ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.src_payload1(\rsp_mux_001|src_payload~93_combout ));

Computer_System_altera_merlin_traffic_limiter_1 arm_a9_hps_h2f_axi_master_wr_limiter(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_WLAST_0(h2f_WLAST_0),
	.clk(outclk_wire_0),
	.Equal0(\router|Equal0~6_combout ),
	.Equal01(\router|Equal0~7_combout ),
	.Equal02(\router|Equal0~14_combout ),
	.sink_ready(\cmd_demux|sink_ready~2_combout ),
	.last_channel_0(\arm_a9_hps_h2f_axi_master_wr_limiter|last_channel[0]~q ),
	.has_pending_responses1(\arm_a9_hps_h2f_axi_master_wr_limiter|has_pending_responses~q ),
	.cmd_sink_ready(\arm_a9_hps_h2f_axi_master_wr_limiter|cmd_sink_ready~0_combout ),
	.out_valid(\onchip_sram_s2_rsp_width_adapter|out_valid~0_combout ),
	.src_payload(\rsp_mux_001|src_payload~0_combout ),
	.src0_valid(\rsp_demux_001|src0_valid~0_combout ),
	.mem_126_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][126]~q ),
	.src0_valid1(\rsp_demux|src0_valid~0_combout ),
	.WideOr1(WideOr1),
	.last_cycle(\cmd_mux|last_cycle~1_combout ),
	.cmd_sink_channel({gnd,\router|Equal0~17_combout }),
	.last_channel_1(\arm_a9_hps_h2f_axi_master_wr_limiter|last_channel[1]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.sink_ready1(\cmd_demux|sink_ready~3_combout ));

Computer_System_Computer_System_mm_interconnect_0_router router(
	.h2f_AWADDR_2(h2f_AWADDR_2),
	.h2f_AWADDR_3(h2f_AWADDR_3),
	.h2f_AWADDR_4(h2f_AWADDR_4),
	.h2f_AWADDR_5(h2f_AWADDR_5),
	.h2f_AWADDR_6(h2f_AWADDR_6),
	.h2f_AWADDR_7(h2f_AWADDR_7),
	.h2f_AWADDR_8(h2f_AWADDR_8),
	.h2f_AWADDR_9(h2f_AWADDR_9),
	.h2f_AWADDR_10(h2f_AWADDR_10),
	.h2f_AWADDR_11(h2f_AWADDR_11),
	.h2f_AWADDR_12(h2f_AWADDR_12),
	.h2f_AWADDR_13(h2f_AWADDR_13),
	.h2f_AWADDR_14(h2f_AWADDR_14),
	.h2f_AWADDR_15(h2f_AWADDR_15),
	.h2f_AWADDR_16(h2f_AWADDR_16),
	.h2f_AWADDR_17(h2f_AWADDR_17),
	.h2f_AWADDR_18(h2f_AWADDR_18),
	.h2f_AWADDR_19(h2f_AWADDR_19),
	.h2f_AWADDR_20(h2f_AWADDR_20),
	.h2f_AWADDR_21(h2f_AWADDR_21),
	.h2f_AWADDR_22(h2f_AWADDR_22),
	.h2f_AWADDR_23(h2f_AWADDR_23),
	.h2f_AWADDR_24(h2f_AWADDR_24),
	.h2f_AWADDR_25(h2f_AWADDR_25),
	.h2f_AWADDR_26(h2f_AWADDR_26),
	.h2f_AWADDR_27(h2f_AWADDR_27),
	.address_burst_24(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[24]~q ),
	.address_burst_25(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[25]~q ),
	.address_burst_23(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[23]~q ),
	.address_burst_13(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[13]~q ),
	.address_burst_21(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[21]~q ),
	.address_burst_22(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[22]~q ),
	.address_burst_19(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[19]~q ),
	.address_burst_20(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[20]~q ),
	.address_burst_15(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[15]~q ),
	.address_burst_16(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[16]~q ),
	.address_burst_17(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[17]~q ),
	.address_burst_18(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[18]~q ),
	.address_burst_26(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[26]~q ),
	.address_burst_27(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[27]~q ),
	.address_burst_12(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[12]~q ),
	.address_burst_14(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[14]~q ),
	.address_burst_10(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[10]~q ),
	.address_burst_11(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[11]~q ),
	.address_burst_9(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[9]~q ),
	.address_burst_8(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[8]~q ),
	.sop_enable(\arm_a9_hps_h2f_axi_master_agent|sop_enable~q ),
	.Equal0(\router|Equal0~6_combout ),
	.Equal01(\router|Equal0~7_combout ),
	.address_burst_7(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[7]~q ),
	.address_burst_6(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[6]~q ),
	.address_burst_2(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[2]~q ),
	.address_burst_3(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[3]~q ),
	.address_burst_4(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[4]~q ),
	.address_burst_5(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[5]~q ),
	.Equal02(\router|Equal0~14_combout ),
	.Equal03(\router|Equal0~16_combout ),
	.Equal04(\router|Equal0~17_combout ));

Computer_System_altera_avalon_sc_fifo_2 onchip_sram_s2_agent_rdata_fifo(
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.clk(outclk_wire_0),
	.read_latency_shift_reg_0(\onchip_sram_s2_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\onchip_sram_s2_agent_rdata_fifo|mem_used[0]~q ),
	.mem_125_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][125]~q ),
	.mem_used_01(\onchip_sram_s2_agent_rsp_fifo|mem_used[0]~q ),
	.out_valid(\onchip_sram_s2_rsp_width_adapter|out_valid~0_combout ),
	.src_payload(\rsp_mux_001|src_payload~0_combout ),
	.always10(\onchip_sram_s2_rsp_width_adapter|always10~9_combout ),
	.always4(\onchip_sram_s2_agent_rdata_fifo|always4~0_combout ),
	.mem_0_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][0]~q ),
	.mem_1_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][1]~q ),
	.mem_2_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][2]~q ),
	.mem_3_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][3]~q ),
	.mem_4_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][4]~q ),
	.mem_5_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][5]~q ),
	.mem_6_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][6]~q ),
	.mem_7_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][7]~q ),
	.mem_8_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][8]~q ),
	.mem_9_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][9]~q ),
	.mem_10_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][10]~q ),
	.mem_11_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][11]~q ),
	.mem_12_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][12]~q ),
	.mem_13_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][13]~q ),
	.mem_14_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][14]~q ),
	.mem_15_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][15]~q ),
	.mem_16_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][16]~q ),
	.mem_17_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][17]~q ),
	.mem_18_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][18]~q ),
	.mem_19_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][19]~q ),
	.mem_20_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][20]~q ),
	.mem_21_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][21]~q ),
	.mem_22_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][22]~q ),
	.mem_23_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][23]~q ),
	.mem_24_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][24]~q ),
	.mem_25_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][25]~q ),
	.mem_26_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][26]~q ),
	.mem_27_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][27]~q ),
	.mem_28_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][28]~q ),
	.mem_29_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][29]~q ),
	.mem_30_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][30]~q ),
	.mem_31_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][31]~q ),
	.out_data_1(\onchip_sram_s2_agent_rdata_fifo|out_data[1]~0_combout ),
	.out_data_4(\onchip_sram_s2_agent_rdata_fifo|out_data[4]~1_combout ),
	.out_data_6(\onchip_sram_s2_agent_rdata_fifo|out_data[6]~2_combout ),
	.out_data_8(\onchip_sram_s2_agent_rdata_fifo|out_data[8]~3_combout ),
	.out_data_13(\onchip_sram_s2_agent_rdata_fifo|out_data[13]~4_combout ),
	.out_data_17(\onchip_sram_s2_agent_rdata_fifo|out_data[17]~5_combout ),
	.out_data_20(\onchip_sram_s2_agent_rdata_fifo|out_data[20]~6_combout ),
	.out_data_22(\onchip_sram_s2_agent_rdata_fifo|out_data[22]~7_combout ),
	.out_data_24(\onchip_sram_s2_agent_rdata_fifo|out_data[24]~8_combout ),
	.out_data_29(\onchip_sram_s2_agent_rdata_fifo|out_data[29]~9_combout ),
	.reset(r_sync_rst),
	.p1_ready(\onchip_sram_s2_rsp_width_adapter|p1_ready~0_combout ));

Computer_System_altera_avalon_sc_fifo_3 onchip_sram_s2_agent_rsp_fifo(
	.clk(outclk_wire_0),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.out_uncomp_byte_cnt_reg_6(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_2(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_3(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_7(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[7]~q ),
	.out_uncomp_byte_cnt_reg_4(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_8(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[8]~q ),
	.out_uncomp_byte_cnt_reg_5(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_burstwrap_reg_2(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[2]~q ),
	.out_burstwrap_reg_3(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[3]~q ),
	.out_addr_reg_1(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[1]~q ),
	.out_burstwrap_reg_1(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[1]~q ),
	.out_addr_reg_0(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[0]~q ),
	.out_burstwrap_reg_0(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[0]~q ),
	.stateST_COMP_TRANS(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.in_data_reg_91(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.in_data_reg_90(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ),
	.mem_used_1(\onchip_sram_s2_agent_rsp_fifo|mem_used[1]~q ),
	.cp_ready(\onchip_sram_s2_agent|cp_ready~combout ),
	.in_eop_reg(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_eop_reg~q ),
	.new_burst_reg(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|new_burst_reg~q ),
	.in_bytecount_reg_zero(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_bytecount_reg_zero~q ),
	.out_valid_reg(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_125_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][125]~q ),
	.mem_used_0(\onchip_sram_s2_agent_rsp_fifo|mem_used[0]~q ),
	.out_valid(\onchip_sram_s2_rsp_width_adapter|out_valid~0_combout ),
	.comb(\onchip_sram_s2_agent|comb~0_combout ),
	.mem_126_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][126]~q ),
	.mem_66_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][66]~q ),
	.mem_80_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][80]~q ),
	.mem_79_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][79]~q ),
	.mem_78_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][74]~q ),
	.mem_38_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][38]~q ),
	.mem_122_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][122]~q ),
	.mem_123_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][123]~q ),
	.mem_91_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][91]~q ),
	.mem_124_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][124]~q ),
	.mem_90_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][90]~q ),
	.mem_39_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][39]~q ),
	.always10(\onchip_sram_s2_rsp_width_adapter|always10~9_combout ),
	.mem_68_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][68]~q ),
	.mem_101_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][101]~q ),
	.mem_102_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][102]~q ),
	.mem_103_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][103]~q ),
	.mem_104_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][104]~q ),
	.mem_105_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][112]~q ),
	.in_data_reg_68(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.reset(r_sync_rst),
	.nxt_out_eop(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~1_combout ),
	.in_data_reg_69(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.last_packet_beat(\onchip_sram_s2_agent|uncompressor|last_packet_beat~5_combout ),
	.p1_ready(\onchip_sram_s2_rsp_width_adapter|p1_ready~0_combout ),
	.cp_ready1(\onchip_sram_s2_agent|cp_ready~0_combout ),
	.out_byte_cnt_reg_2(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.WideOr0(\onchip_sram_s2_agent|WideOr0~combout ),
	.always101(\onchip_sram_s2_rsp_width_adapter|always10~10_combout ),
	.mem_83_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][83]~q ),
	.in_data_reg_122(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[122]~q ),
	.in_data_reg_123(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[123]~q ),
	.in_data_reg_124(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[124]~q ),
	.mem_84_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][84]~q ),
	.in_data_reg_101(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.in_data_reg_104(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[104]~q ),
	.in_data_reg_105(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.mem_37_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][37]~q ),
	.mem_82_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][82]~q ),
	.mem_36_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][36]~q ),
	.mem_81_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][81]~q ));

Computer_System_altera_merlin_slave_agent_1 onchip_sram_s2_agent(
	.outclk_wire_0(outclk_wire_0),
	.in_ready_hold(in_ready_hold),
	.in_narrow_reg(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.always12(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|always12~0_combout ),
	.in_byteen_reg_2(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.source0_data_34(source0_data_34),
	.in_byteen_reg_0(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.source0_data_32(source0_data_32),
	.in_byteen_reg_1(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.source0_data_33(source0_data_33),
	.in_byteen_reg_3(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.source0_data_35(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~3_combout ),
	.source0_data_351(source0_data_35),
	.mem_used_1(\onchip_sram_s2_agent_rsp_fifo|mem_used[1]~q ),
	.cp_ready1(\onchip_sram_s2_agent|cp_ready~combout ),
	.out_valid_reg(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.ShiftLeft1(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|ShiftLeft1~0_combout ),
	.source0_data_352(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|source0_data[35]~5_combout ),
	.WideOr01(\onchip_sram_s2_agent|WideOr0~0_combout ),
	.read_latency_shift_reg_0(\onchip_sram_s2_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\onchip_sram_s2_agent_rdata_fifo|mem_used[0]~q ),
	.mem_125_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][125]~q ),
	.mem_used_01(\onchip_sram_s2_agent_rsp_fifo|mem_used[0]~q ),
	.out_valid(\onchip_sram_s2_rsp_width_adapter|out_valid~0_combout ),
	.comb(\onchip_sram_s2_agent|comb~0_combout ),
	.mem_66_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][66]~q ),
	.burst_uncompress_busy(\onchip_sram_s2_agent|uncompressor|burst_uncompress_busy~q ),
	.last_packet_beat(\onchip_sram_s2_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat1(\onchip_sram_s2_agent|uncompressor|last_packet_beat~1_combout ),
	.mem_80_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][80]~q ),
	.mem_79_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][79]~q ),
	.mem_78_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][78]~q ),
	.mem_77_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][77]~q ),
	.mem_76_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][76]~q ),
	.mem_75_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][75]~q ),
	.mem_74_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][74]~q ),
	.last_packet_beat2(\onchip_sram_s2_agent|uncompressor|last_packet_beat~4_combout ),
	.src_payload(\rsp_mux_001|src_payload~0_combout ),
	.mem_38_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][38]~q ),
	.source_addr_2(\onchip_sram_s2_agent|uncompressor|source_addr[2]~0_combout ),
	.source_addr_21(\onchip_sram_s2_agent|uncompressor|source_addr[2]~1_combout ),
	.mem_91_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][91]~q ),
	.mem_90_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][90]~q ),
	.mem_39_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][39]~q ),
	.source_addr_3(\onchip_sram_s2_agent|uncompressor|source_addr[3]~2_combout ),
	.always10(\onchip_sram_s2_rsp_width_adapter|always10~9_combout ),
	.in_data_reg_68(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.m0_write(m0_write1),
	.r_sync_rst(r_sync_rst),
	.last_packet_beat3(\onchip_sram_s2_agent|uncompressor|last_packet_beat~5_combout ),
	.p1_ready(\onchip_sram_s2_rsp_width_adapter|p1_ready~0_combout ),
	.cp_ready2(\onchip_sram_s2_agent|cp_ready~0_combout ),
	.cp_ready3(\onchip_sram_s2_agent|cp_ready~1_combout ),
	.WideOr02(\onchip_sram_s2_agent|WideOr0~combout ),
	.mem_83_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][83]~q ),
	.mem_84_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][84]~q ),
	.mem_37_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][37]~q ),
	.mem_82_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][82]~q ),
	.mem_36_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][36]~q ),
	.mem_81_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][81]~q ));

Computer_System_altera_avalon_sc_fifo fifo_hps_to_fpga_in_agent_rdata_fifo(
	.clk(outclk_wire_0),
	.in_ready_hold(in_ready_hold),
	.mem_31_0(\fifo_hps_to_fpga_in_agent_rdata_fifo|mem[0][31]~q ),
	.reset(r_sync_rst));

Computer_System_altera_avalon_sc_fifo_1 fifo_hps_to_fpga_in_agent_rsp_fifo(
	.clk(outclk_wire_0),
	.out_valid_reg(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem_used[1]~q ),
	.mem_68_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][68]~q ),
	.mem_125_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][125]~q ),
	.mem_used_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem_used[0]~q ),
	.comb(\fifo_hps_to_fpga_in_agent|comb~0_combout ),
	.mem_122_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][122]~q ),
	.mem_123_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][123]~q ),
	.mem_124_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][124]~q ),
	.mem_90_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][90]~q ),
	.mem_91_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][91]~q ),
	.ShiftRight0(\fifo_hps_to_fpga_in_rsp_width_adapter|ShiftRight0~0_combout ),
	.mem_38_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][38]~q ),
	.always10(\fifo_hps_to_fpga_in_rsp_width_adapter|always10~0_combout ),
	.mem_126_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][126]~q ),
	.mem_39_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][39]~q ),
	.always101(\fifo_hps_to_fpga_in_rsp_width_adapter|always10~1_combout ),
	.mem_101_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][101]~q ),
	.mem_102_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][102]~q ),
	.mem_103_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][103]~q ),
	.mem_104_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][104]~q ),
	.mem_105_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][112]~q ),
	.in_data_reg_68(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.nxt_uncomp_subburst_byte_cnt(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_uncomp_subburst_byte_cnt~0_combout ),
	.reset(r_sync_rst),
	.in_eop_reg(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_eop_reg~q ),
	.cp_ready(\fifo_hps_to_fpga_in_agent|cp_ready~0_combout ),
	.p1_ready(\fifo_hps_to_fpga_in_rsp_width_adapter|p1_ready~0_combout ),
	.read(\fifo_hps_to_fpga_in_agent_rsp_fifo|read~0_combout ),
	.always102(\fifo_hps_to_fpga_in_rsp_width_adapter|always10~2_combout ),
	.in_data_reg_122(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[122]~q ),
	.in_data_reg_123(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[123]~q ),
	.in_data_reg_124(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[124]~q ),
	.in_data_reg_90(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ),
	.in_data_reg_91(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.int_nxt_addr_reg_dly_2(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.mem_83_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][83]~q ),
	.int_nxt_addr_reg_dly_3(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.mem_84_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][84]~q ),
	.in_data_reg_101(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.in_data_reg_104(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[104]~q ),
	.in_data_reg_105(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[105]~q ),
	.in_data_reg_106(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[106]~q ),
	.in_data_reg_107(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[107]~q ),
	.in_data_reg_108(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[108]~q ),
	.in_data_reg_109(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[109]~q ),
	.in_data_reg_110(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[110]~q ),
	.in_data_reg_111(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[111]~q ),
	.in_data_reg_112(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[112]~q ),
	.out_burstwrap_reg_2(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[2]~q ),
	.out_burstwrap_reg_3(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[3]~q ),
	.mem_37_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][37]~q ),
	.out_addr_reg_1(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[1]~q ),
	.mem_82_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][82]~q ),
	.mem_36_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][36]~q ),
	.out_burstwrap_reg_1(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[1]~q ),
	.out_addr_reg_0(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_addr_reg[0]~q ),
	.mem_81_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][81]~q ),
	.out_burstwrap_reg_0(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_burstwrap_reg[0]~q ));

Computer_System_altera_merlin_slave_agent fifo_hps_to_fpga_in_agent(
	.outclk_wire_0(outclk_wire_0),
	.op_2(op_2),
	.op_21(op_21),
	.op_22(op_22),
	.in_byteen_reg_3(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\fifo_hps_to_fpga_in_agent|WideOr0~0_combout ),
	.wrfull(wrfull),
	.wrfull1(wrfull2),
	.mem_used_1(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem_used[1]~q ),
	.mem_125_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][125]~q ),
	.mem_used_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem_used[0]~q ),
	.comb(\fifo_hps_to_fpga_in_agent|comb~0_combout ),
	.mem_90_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][90]~q ),
	.mem_91_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][91]~q ),
	.mem_38_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][38]~q ),
	.source_addr_2(\fifo_hps_to_fpga_in_agent|uncompressor|source_addr[2]~0_combout ),
	.mem_39_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][39]~q ),
	.source_addr_3(\fifo_hps_to_fpga_in_agent|uncompressor|source_addr[3]~1_combout ),
	.in_data_reg_68(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[68]~q ),
	.nxt_uncomp_subburst_byte_cnt(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_uncomp_subburst_byte_cnt~0_combout ),
	.m0_write(m0_write),
	.r_sync_rst(r_sync_rst),
	.wrfull2(wrfull4),
	.cp_ready(\fifo_hps_to_fpga_in_agent|cp_ready~0_combout ),
	.read(\fifo_hps_to_fpga_in_agent_rsp_fifo|read~0_combout ),
	.cp_ready1(\fifo_hps_to_fpga_in_agent|cp_ready~1_combout ),
	.mem_83_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][83]~q ),
	.mem_84_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][84]~q ),
	.mem_37_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][37]~q ),
	.mem_82_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][82]~q ),
	.mem_36_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][36]~q ),
	.mem_81_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][81]~q ));

Computer_System_altera_merlin_axi_master_ni arm_a9_hps_h2f_axi_master_agent(
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_ARLEN_0(h2f_ARLEN_0),
	.h2f_ARLEN_1(h2f_ARLEN_1),
	.h2f_ARLEN_2(h2f_ARLEN_2),
	.h2f_ARLEN_3(h2f_ARLEN_3),
	.h2f_ARSIZE_0(h2f_ARSIZE_0),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWADDR_0(h2f_AWADDR_0),
	.h2f_AWADDR_1(h2f_AWADDR_1),
	.h2f_AWADDR_2(h2f_AWADDR_2),
	.h2f_AWADDR_3(h2f_AWADDR_3),
	.h2f_AWADDR_4(h2f_AWADDR_4),
	.h2f_AWADDR_5(h2f_AWADDR_5),
	.h2f_AWADDR_6(h2f_AWADDR_6),
	.h2f_AWADDR_7(h2f_AWADDR_7),
	.h2f_AWADDR_8(h2f_AWADDR_8),
	.h2f_AWADDR_9(h2f_AWADDR_9),
	.h2f_AWADDR_10(h2f_AWADDR_10),
	.h2f_AWADDR_11(h2f_AWADDR_11),
	.h2f_AWADDR_12(h2f_AWADDR_12),
	.h2f_AWADDR_13(h2f_AWADDR_13),
	.h2f_AWADDR_14(h2f_AWADDR_14),
	.h2f_AWADDR_15(h2f_AWADDR_15),
	.h2f_AWADDR_16(h2f_AWADDR_16),
	.h2f_AWADDR_17(h2f_AWADDR_17),
	.h2f_AWADDR_18(h2f_AWADDR_18),
	.h2f_AWADDR_19(h2f_AWADDR_19),
	.h2f_AWADDR_20(h2f_AWADDR_20),
	.h2f_AWADDR_21(h2f_AWADDR_21),
	.h2f_AWADDR_22(h2f_AWADDR_22),
	.h2f_AWADDR_23(h2f_AWADDR_23),
	.h2f_AWADDR_24(h2f_AWADDR_24),
	.h2f_AWADDR_25(h2f_AWADDR_25),
	.h2f_AWADDR_26(h2f_AWADDR_26),
	.h2f_AWADDR_27(h2f_AWADDR_27),
	.h2f_AWBURST_0(h2f_AWBURST_0),
	.h2f_AWBURST_1(h2f_AWBURST_1),
	.h2f_AWLEN_0(h2f_AWLEN_0),
	.h2f_AWLEN_1(h2f_AWLEN_1),
	.h2f_AWLEN_2(h2f_AWLEN_2),
	.h2f_AWLEN_3(h2f_AWLEN_3),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.outclk_wire_0(outclk_wire_0),
	.address_burst_24(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[24]~q ),
	.address_burst_25(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[25]~q ),
	.address_burst_23(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[23]~q ),
	.address_burst_13(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[13]~q ),
	.address_burst_21(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[21]~q ),
	.address_burst_22(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[22]~q ),
	.address_burst_19(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[19]~q ),
	.address_burst_20(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[20]~q ),
	.address_burst_15(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[15]~q ),
	.address_burst_16(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[16]~q ),
	.address_burst_17(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[17]~q ),
	.address_burst_18(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[18]~q ),
	.address_burst_26(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[26]~q ),
	.address_burst_27(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[27]~q ),
	.address_burst_12(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[12]~q ),
	.address_burst_14(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[14]~q ),
	.address_burst_10(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[10]~q ),
	.address_burst_11(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[11]~q ),
	.address_burst_9(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[9]~q ),
	.address_burst_8(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[8]~q ),
	.Add4(\arm_a9_hps_h2f_axi_master_agent|Add4~1_sumout ),
	.Add5(\arm_a9_hps_h2f_axi_master_agent|Add5~1_sumout ),
	.Add41(\arm_a9_hps_h2f_axi_master_agent|Add4~5_sumout ),
	.Add51(\arm_a9_hps_h2f_axi_master_agent|Add5~5_sumout ),
	.Add42(\arm_a9_hps_h2f_axi_master_agent|Add4~9_sumout ),
	.Add52(\arm_a9_hps_h2f_axi_master_agent|Add5~9_sumout ),
	.Add43(\arm_a9_hps_h2f_axi_master_agent|Add4~13_sumout ),
	.Add53(\arm_a9_hps_h2f_axi_master_agent|Add5~13_sumout ),
	.Add44(\arm_a9_hps_h2f_axi_master_agent|Add4~17_sumout ),
	.Add54(\arm_a9_hps_h2f_axi_master_agent|Add5~17_sumout ),
	.Add55(\arm_a9_hps_h2f_axi_master_agent|Add5~21_sumout ),
	.Add45(\arm_a9_hps_h2f_axi_master_agent|Add4~21_sumout ),
	.Add56(\arm_a9_hps_h2f_axi_master_agent|Add5~25_sumout ),
	.Add46(\arm_a9_hps_h2f_axi_master_agent|Add4~25_sumout ),
	.Add47(\arm_a9_hps_h2f_axi_master_agent|Add4~29_sumout ),
	.Add57(\arm_a9_hps_h2f_axi_master_agent|Add5~29_sumout ),
	.Add48(\arm_a9_hps_h2f_axi_master_agent|Add4~33_sumout ),
	.Add58(\arm_a9_hps_h2f_axi_master_agent|Add5~33_sumout ),
	.in_ready(\onchip_sram_s2_cmd_width_adapter|in_ready~0_combout ),
	.nxt_in_ready(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~4_combout ),
	.sop_enable1(\arm_a9_hps_h2f_axi_master_agent|sop_enable~q ),
	.address_burst_7(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[7]~q ),
	.address_burst_6(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[6]~q ),
	.address_burst_2(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[2]~q ),
	.address_burst_3(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[3]~q ),
	.address_burst_4(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[4]~q ),
	.address_burst_5(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[5]~q ),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.sink_ready1(\cmd_demux|sink_ready~2_combout ),
	.cmd_sink_ready(\arm_a9_hps_h2f_axi_master_wr_limiter|cmd_sink_ready~0_combout ),
	.last_cycle(\cmd_mux|last_cycle~0_combout ),
	.awready(ARM_A9_HPS_h2f_axi_master_awready),
	.last_cycle1(\cmd_mux|last_cycle~1_combout ),
	.wready(ARM_A9_HPS_h2f_axi_master_wready),
	.LessThan11(\arm_a9_hps_h2f_axi_master_agent|LessThan11~0_combout ),
	.Add3(\arm_a9_hps_h2f_axi_master_agent|Add3~0_combout ),
	.log2ceil(\arm_a9_hps_h2f_axi_master_agent|log2ceil~0_combout ),
	.address_burst_1(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[1]~q ),
	.LessThan10(\arm_a9_hps_h2f_axi_master_agent|LessThan10~0_combout ),
	.Add31(\arm_a9_hps_h2f_axi_master_agent|Add3~1_combout ),
	.address_burst_0(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[0]~q ),
	.out_data_2(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[2]~0_combout ),
	.out_data_3(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[3]~1_combout ),
	.burst_bytecount_4(\arm_a9_hps_h2f_axi_master_agent|burst_bytecount[4]~q ),
	.burst_bytecount_6(\arm_a9_hps_h2f_axi_master_agent|burst_bytecount[6]~q ),
	.burst_bytecount_5(\arm_a9_hps_h2f_axi_master_agent|burst_bytecount[5]~q ),
	.burst_bytecount_7(\arm_a9_hps_h2f_axi_master_agent|burst_bytecount[7]~q ),
	.Add0(\arm_a9_hps_h2f_axi_master_agent|Add0~0_combout ),
	.Add2(\arm_a9_hps_h2f_axi_master_agent|Add2~0_combout ),
	.Add01(\arm_a9_hps_h2f_axi_master_agent|Add0~1_combout ),
	.Add21(\arm_a9_hps_h2f_axi_master_agent|Add2~1_combout ),
	.Add22(\arm_a9_hps_h2f_axi_master_agent|Add2~2_combout ),
	.write_cp_data_188(\arm_a9_hps_h2f_axi_master_agent|write_cp_data[188]~0_combout ),
	.write_cp_data_187(\arm_a9_hps_h2f_axi_master_agent|write_cp_data[187]~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.out_data_7(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[7]~20_combout ),
	.Add1(\arm_a9_hps_h2f_axi_master_agent|Add1~3_combout ),
	.out_data_9(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[9]~21_combout ),
	.out_data_6(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[6]~22_combout ),
	.LessThan16(\arm_a9_hps_h2f_axi_master_agent|LessThan16~0_combout ),
	.out_data_8(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[8]~23_combout ),
	.LessThan12(\arm_a9_hps_h2f_axi_master_agent|LessThan12~0_combout ),
	.Selector26(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|Selector26~0_combout ),
	.out_data_4(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[4]~24_combout ),
	.LessThan14(\arm_a9_hps_h2f_axi_master_agent|LessThan14~0_combout ),
	.out_data_5(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[5]~25_combout ),
	.LessThan15(\arm_a9_hps_h2f_axi_master_agent|LessThan15~0_combout ),
	.LessThan2(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|LessThan2~0_combout ),
	.Add32(\arm_a9_hps_h2f_axi_master_agent|Add3~2_combout ),
	.Selector7(\arm_a9_hps_h2f_axi_master_agent|Selector7~0_combout ),
	.out_data_1(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[1]~26_combout ),
	.Decoder0(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|Decoder0~1_combout ),
	.Selector8(\arm_a9_hps_h2f_axi_master_agent|Selector8~0_combout ),
	.out_data_0(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[0]~27_combout ),
	.Selector6(\arm_a9_hps_h2f_axi_master_agent|Selector6~0_combout ),
	.Selector5(\arm_a9_hps_h2f_axi_master_agent|Selector5~0_combout ));

Computer_System_altera_merlin_slave_translator_1 onchip_sram_s2_translator(
	.clk(outclk_wire_0),
	.in_ready_hold(in_ready_hold),
	.mem_used_1(\onchip_sram_s2_agent_rsp_fifo|mem_used[1]~q ),
	.out_valid_reg(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.read_latency_shift_reg_0(\onchip_sram_s2_translator|read_latency_shift_reg[0]~q ),
	.reset(r_sync_rst),
	.in_data_reg_69(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[69]~q ),
	.WideOr0(\onchip_sram_s2_agent|WideOr0~combout ));

Computer_System_altera_merlin_width_adapter_2 onchip_sram_s2_cmd_width_adapter(
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_ARADDR_1(h2f_ARADDR_1),
	.h2f_ARADDR_3(h2f_ARADDR_3),
	.h2f_ARSIZE_1(h2f_ARSIZE_1),
	.h2f_ARSIZE_2(h2f_ARSIZE_2),
	.h2f_AWADDR_1(h2f_AWADDR_1),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.h2f_WDATA_0(h2f_WDATA_0),
	.h2f_WDATA_1(h2f_WDATA_1),
	.h2f_WDATA_2(h2f_WDATA_2),
	.h2f_WDATA_3(h2f_WDATA_3),
	.h2f_WDATA_4(h2f_WDATA_4),
	.h2f_WDATA_5(h2f_WDATA_5),
	.h2f_WDATA_6(h2f_WDATA_6),
	.h2f_WDATA_7(h2f_WDATA_7),
	.h2f_WDATA_8(h2f_WDATA_8),
	.h2f_WDATA_9(h2f_WDATA_9),
	.h2f_WDATA_10(h2f_WDATA_10),
	.h2f_WDATA_11(h2f_WDATA_11),
	.h2f_WDATA_12(h2f_WDATA_12),
	.h2f_WDATA_13(h2f_WDATA_13),
	.h2f_WDATA_14(h2f_WDATA_14),
	.h2f_WDATA_15(h2f_WDATA_15),
	.h2f_WDATA_16(h2f_WDATA_16),
	.h2f_WDATA_17(h2f_WDATA_17),
	.h2f_WDATA_18(h2f_WDATA_18),
	.h2f_WDATA_19(h2f_WDATA_19),
	.h2f_WDATA_20(h2f_WDATA_20),
	.h2f_WDATA_21(h2f_WDATA_21),
	.h2f_WDATA_22(h2f_WDATA_22),
	.h2f_WDATA_23(h2f_WDATA_23),
	.h2f_WDATA_24(h2f_WDATA_24),
	.h2f_WDATA_25(h2f_WDATA_25),
	.h2f_WDATA_26(h2f_WDATA_26),
	.h2f_WDATA_27(h2f_WDATA_27),
	.h2f_WDATA_28(h2f_WDATA_28),
	.h2f_WDATA_29(h2f_WDATA_29),
	.h2f_WDATA_30(h2f_WDATA_30),
	.h2f_WDATA_31(h2f_WDATA_31),
	.h2f_WDATA_32(h2f_WDATA_32),
	.h2f_WDATA_33(h2f_WDATA_33),
	.h2f_WDATA_34(h2f_WDATA_34),
	.h2f_WDATA_35(h2f_WDATA_35),
	.h2f_WDATA_36(h2f_WDATA_36),
	.h2f_WDATA_37(h2f_WDATA_37),
	.h2f_WDATA_38(h2f_WDATA_38),
	.h2f_WDATA_39(h2f_WDATA_39),
	.h2f_WDATA_40(h2f_WDATA_40),
	.h2f_WDATA_41(h2f_WDATA_41),
	.h2f_WDATA_42(h2f_WDATA_42),
	.h2f_WDATA_43(h2f_WDATA_43),
	.h2f_WDATA_44(h2f_WDATA_44),
	.h2f_WDATA_45(h2f_WDATA_45),
	.h2f_WDATA_46(h2f_WDATA_46),
	.h2f_WDATA_47(h2f_WDATA_47),
	.h2f_WDATA_48(h2f_WDATA_48),
	.h2f_WDATA_49(h2f_WDATA_49),
	.h2f_WDATA_50(h2f_WDATA_50),
	.h2f_WDATA_51(h2f_WDATA_51),
	.h2f_WDATA_52(h2f_WDATA_52),
	.h2f_WDATA_53(h2f_WDATA_53),
	.h2f_WDATA_54(h2f_WDATA_54),
	.h2f_WDATA_55(h2f_WDATA_55),
	.h2f_WDATA_56(h2f_WDATA_56),
	.h2f_WDATA_57(h2f_WDATA_57),
	.h2f_WDATA_58(h2f_WDATA_58),
	.h2f_WDATA_59(h2f_WDATA_59),
	.h2f_WDATA_60(h2f_WDATA_60),
	.h2f_WDATA_61(h2f_WDATA_61),
	.h2f_WDATA_62(h2f_WDATA_62),
	.h2f_WDATA_63(h2f_WDATA_63),
	.h2f_WDATA_64(h2f_WDATA_64),
	.h2f_WDATA_65(h2f_WDATA_65),
	.h2f_WDATA_66(h2f_WDATA_66),
	.h2f_WDATA_67(h2f_WDATA_67),
	.h2f_WDATA_68(h2f_WDATA_68),
	.h2f_WDATA_69(h2f_WDATA_69),
	.h2f_WDATA_70(h2f_WDATA_70),
	.h2f_WDATA_71(h2f_WDATA_71),
	.h2f_WDATA_72(h2f_WDATA_72),
	.h2f_WDATA_73(h2f_WDATA_73),
	.h2f_WDATA_74(h2f_WDATA_74),
	.h2f_WDATA_75(h2f_WDATA_75),
	.h2f_WDATA_76(h2f_WDATA_76),
	.h2f_WDATA_77(h2f_WDATA_77),
	.h2f_WDATA_78(h2f_WDATA_78),
	.h2f_WDATA_79(h2f_WDATA_79),
	.h2f_WDATA_80(h2f_WDATA_80),
	.h2f_WDATA_81(h2f_WDATA_81),
	.h2f_WDATA_82(h2f_WDATA_82),
	.h2f_WDATA_83(h2f_WDATA_83),
	.h2f_WDATA_84(h2f_WDATA_84),
	.h2f_WDATA_85(h2f_WDATA_85),
	.h2f_WDATA_86(h2f_WDATA_86),
	.h2f_WDATA_87(h2f_WDATA_87),
	.h2f_WDATA_88(h2f_WDATA_88),
	.h2f_WDATA_89(h2f_WDATA_89),
	.h2f_WDATA_90(h2f_WDATA_90),
	.h2f_WDATA_91(h2f_WDATA_91),
	.h2f_WDATA_92(h2f_WDATA_92),
	.h2f_WDATA_93(h2f_WDATA_93),
	.h2f_WDATA_94(h2f_WDATA_94),
	.h2f_WDATA_95(h2f_WDATA_95),
	.h2f_WDATA_96(h2f_WDATA_96),
	.h2f_WDATA_97(h2f_WDATA_97),
	.h2f_WDATA_98(h2f_WDATA_98),
	.h2f_WDATA_99(h2f_WDATA_99),
	.h2f_WDATA_100(h2f_WDATA_100),
	.h2f_WDATA_101(h2f_WDATA_101),
	.h2f_WDATA_102(h2f_WDATA_102),
	.h2f_WDATA_103(h2f_WDATA_103),
	.h2f_WDATA_104(h2f_WDATA_104),
	.h2f_WDATA_105(h2f_WDATA_105),
	.h2f_WDATA_106(h2f_WDATA_106),
	.h2f_WDATA_107(h2f_WDATA_107),
	.h2f_WDATA_108(h2f_WDATA_108),
	.h2f_WDATA_109(h2f_WDATA_109),
	.h2f_WDATA_110(h2f_WDATA_110),
	.h2f_WDATA_111(h2f_WDATA_111),
	.h2f_WDATA_112(h2f_WDATA_112),
	.h2f_WDATA_113(h2f_WDATA_113),
	.h2f_WDATA_114(h2f_WDATA_114),
	.h2f_WDATA_115(h2f_WDATA_115),
	.h2f_WDATA_116(h2f_WDATA_116),
	.h2f_WDATA_117(h2f_WDATA_117),
	.h2f_WDATA_118(h2f_WDATA_118),
	.h2f_WDATA_119(h2f_WDATA_119),
	.h2f_WDATA_120(h2f_WDATA_120),
	.h2f_WDATA_121(h2f_WDATA_121),
	.h2f_WDATA_122(h2f_WDATA_122),
	.h2f_WDATA_123(h2f_WDATA_123),
	.h2f_WDATA_124(h2f_WDATA_124),
	.h2f_WDATA_125(h2f_WDATA_125),
	.h2f_WDATA_126(h2f_WDATA_126),
	.h2f_WDATA_127(h2f_WDATA_127),
	.outclk_wire_0(outclk_wire_0),
	.Mux4(\onchip_sram_s2_cmd_width_adapter|Mux4~0_combout ),
	.Mux5(\onchip_sram_s2_cmd_width_adapter|Mux5~0_combout ),
	.Mux6(\onchip_sram_s2_cmd_width_adapter|Mux6~0_combout ),
	.Mux7(\onchip_sram_s2_cmd_width_adapter|Mux7~0_combout ),
	.Mux8(\onchip_sram_s2_cmd_width_adapter|Mux8~0_combout ),
	.Mux9(\onchip_sram_s2_cmd_width_adapter|Mux9~0_combout ),
	.Mux10(\onchip_sram_s2_cmd_width_adapter|Mux10~0_combout ),
	.Mux11(\onchip_sram_s2_cmd_width_adapter|Mux11~0_combout ),
	.Mux12(\onchip_sram_s2_cmd_width_adapter|Mux12~0_combout ),
	.Mux13(\onchip_sram_s2_cmd_width_adapter|Mux13~0_combout ),
	.Mux14(\onchip_sram_s2_cmd_width_adapter|Mux14~0_combout ),
	.Mux15(\onchip_sram_s2_cmd_width_adapter|Mux15~0_combout ),
	.Mux16(\onchip_sram_s2_cmd_width_adapter|Mux16~0_combout ),
	.Mux17(\onchip_sram_s2_cmd_width_adapter|Mux17~0_combout ),
	.Mux18(\onchip_sram_s2_cmd_width_adapter|Mux18~0_combout ),
	.Mux19(\onchip_sram_s2_cmd_width_adapter|Mux19~0_combout ),
	.Mux20(\onchip_sram_s2_cmd_width_adapter|Mux20~0_combout ),
	.Mux21(\onchip_sram_s2_cmd_width_adapter|Mux21~0_combout ),
	.Mux22(\onchip_sram_s2_cmd_width_adapter|Mux22~0_combout ),
	.Mux23(\onchip_sram_s2_cmd_width_adapter|Mux23~0_combout ),
	.Mux24(\onchip_sram_s2_cmd_width_adapter|Mux24~0_combout ),
	.Mux25(\onchip_sram_s2_cmd_width_adapter|Mux25~0_combout ),
	.Mux26(\onchip_sram_s2_cmd_width_adapter|Mux26~0_combout ),
	.Mux27(\onchip_sram_s2_cmd_width_adapter|Mux27~0_combout ),
	.Mux28(\onchip_sram_s2_cmd_width_adapter|Mux28~0_combout ),
	.Mux29(\onchip_sram_s2_cmd_width_adapter|Mux29~0_combout ),
	.Mux30(\onchip_sram_s2_cmd_width_adapter|Mux30~0_combout ),
	.Mux31(\onchip_sram_s2_cmd_width_adapter|Mux31~0_combout ),
	.Mux32(\onchip_sram_s2_cmd_width_adapter|Mux32~0_combout ),
	.Mux33(\onchip_sram_s2_cmd_width_adapter|Mux33~0_combout ),
	.Mux34(\onchip_sram_s2_cmd_width_adapter|Mux34~0_combout ),
	.Mux35(\onchip_sram_s2_cmd_width_adapter|Mux35~0_combout ),
	.src_data_185(\cmd_mux_001|src_data[185]~43_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.saved_grant_0(\cmd_mux_001|saved_grant[0]~q ),
	.src_data_198(\cmd_mux_001|src_data[198]~combout ),
	.src_data_199(\cmd_mux_001|src_data[199]~combout ),
	.src_data_200(\cmd_mux_001|src_data[200]~combout ),
	.in_ready(\onchip_sram_s2_cmd_width_adapter|in_ready~0_combout ),
	.nxt_in_ready(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready1(\onchip_sram_s2_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.sop_enable(\arm_a9_hps_h2f_axi_master_agent|sop_enable~q ),
	.r_sync_rst(r_sync_rst),
	.WideOr1(\cmd_mux_001|WideOr1~combout ),
	.in_endofpacket(\cmd_mux_001|src_payload[0]~combout ),
	.use_reg1(\onchip_sram_s2_cmd_width_adapter|use_reg~q ),
	.out_data_91(\onchip_sram_s2_cmd_width_adapter|out_data[91]~0_combout ),
	.out_data_90(\onchip_sram_s2_cmd_width_adapter|out_data[90]~1_combout ),
	.address_burst_1(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|address_burst[1]~q ),
	.out_data_37(\onchip_sram_s2_cmd_width_adapter|out_data[37]~3_combout ),
	.src_data_144(\cmd_mux_001|src_data[144]~combout ),
	.out_data_36(\onchip_sram_s2_cmd_width_adapter|out_data[36]~4_combout ),
	.src_data_130(\cmd_mux_001|src_data[130]~combout ),
	.src_data_134(\cmd_mux_001|src_data[134]~combout ),
	.src_data_138(\cmd_mux_001|src_data[138]~combout ),
	.src_data_142(\cmd_mux_001|src_data[142]~combout ),
	.src_data_146(\cmd_mux_001|src_data[146]~combout ),
	.int_output_sel_0(\onchip_sram_s2_cmd_width_adapter|int_output_sel[0]~0_combout ),
	.out_data_3(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[3]~1_combout ),
	.Mux1(\onchip_sram_s2_cmd_width_adapter|Mux1~0_combout ),
	.src_data_128(\cmd_mux_001|src_data[128]~combout ),
	.src_data_132(\cmd_mux_001|src_data[132]~combout ),
	.src_data_136(\cmd_mux_001|src_data[136]~combout ),
	.src_data_140(\cmd_mux_001|src_data[140]~combout ),
	.Mux3(\onchip_sram_s2_cmd_width_adapter|Mux3~0_combout ),
	.src_data_129(\cmd_mux_001|src_data[129]~combout ),
	.src_data_133(\cmd_mux_001|src_data[133]~combout ),
	.src_data_137(\cmd_mux_001|src_data[137]~combout ),
	.src_data_141(\cmd_mux_001|src_data[141]~combout ),
	.Mux2(\onchip_sram_s2_cmd_width_adapter|Mux2~0_combout ),
	.src_data_131(\cmd_mux_001|src_data[131]~combout ),
	.src_data_135(\cmd_mux_001|src_data[135]~combout ),
	.src_data_139(\cmd_mux_001|src_data[139]~combout ),
	.src_data_143(\cmd_mux_001|src_data[143]~combout ),
	.Mux0(\onchip_sram_s2_cmd_width_adapter|Mux0~0_combout ),
	.out_endofpacket(\onchip_sram_s2_cmd_width_adapter|out_endofpacket~2_combout ),
	.src_data_184(\cmd_mux_001|src_data[184]~combout ),
	.src_payload(\cmd_mux_001|src_payload~2_combout ),
	.src_payload1(\cmd_mux_001|src_payload~3_combout ),
	.src_payload2(\cmd_mux_001|src_payload~4_combout ),
	.src_payload3(\cmd_mux_001|src_payload~5_combout ),
	.out_data_74(\onchip_sram_s2_cmd_width_adapter|out_data[74]~5_combout ),
	.src_data_187(\cmd_mux_001|src_data[187]~combout ),
	.src_data_186(\cmd_mux_001|src_data[186]~combout ),
	.write_cp_data_188(\arm_a9_hps_h2f_axi_master_agent|write_cp_data[188]~0_combout ),
	.src_payload4(\cmd_mux_001|src_payload~6_combout ),
	.src_data_188(\cmd_mux_001|src_data[188]~combout ),
	.out_data_79(\onchip_sram_s2_cmd_width_adapter|out_data[79]~6_combout ),
	.out_data_76(\onchip_sram_s2_cmd_width_adapter|out_data[76]~7_combout ),
	.write_cp_data_187(\arm_a9_hps_h2f_axi_master_agent|write_cp_data[187]~1_combout ),
	.src_payload5(\cmd_mux_001|src_payload~7_combout ),
	.out_data_77(\onchip_sram_s2_cmd_width_adapter|out_data[77]~11_combout ),
	.out_data_78(\onchip_sram_s2_cmd_width_adapter|out_data[78]~14_combout ),
	.out_data_80(\onchip_sram_s2_cmd_width_adapter|out_data[80]~15_combout ),
	.out_data_75(\onchip_sram_s2_cmd_width_adapter|out_data[75]~16_combout ),
	.out_data_7(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[7]~20_combout ),
	.out_data_6(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[6]~22_combout ),
	.out_data_4(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[4]~24_combout ),
	.out_data_5(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[5]~25_combout ),
	.address_reg_4(\onchip_sram_s2_cmd_width_adapter|address_reg[4]~q ),
	.src_payload6(\cmd_mux_001|src_payload~10_combout ),
	.address_reg_5(\onchip_sram_s2_cmd_width_adapter|address_reg[5]~q ),
	.src_payload7(\cmd_mux_001|src_payload~11_combout ),
	.address_reg_6(\onchip_sram_s2_cmd_width_adapter|address_reg[6]~q ),
	.src_payload8(\cmd_mux_001|src_payload~12_combout ),
	.address_reg_7(\onchip_sram_s2_cmd_width_adapter|address_reg[7]~q ),
	.src_payload9(\cmd_mux_001|src_payload~13_combout ),
	.src_data_152(\cmd_mux_001|src_data[152]~combout ),
	.out_data_44(\onchip_sram_s2_cmd_width_adapter|out_data[44]~17_combout ),
	.src_payload10(\cmd_mux_001|src_payload~14_combout ),
	.src_payload11(\cmd_mux_001|src_payload~15_combout ),
	.out_data_45(\onchip_sram_s2_cmd_width_adapter|out_data[45]~18_combout ),
	.int_output_sel_1(\onchip_sram_s2_cmd_width_adapter|int_output_sel[1]~2_combout ));

Computer_System_altera_merlin_width_adapter fifo_hps_to_fpga_in_cmd_width_adapter(
	.h2f_WLAST_0(h2f_WLAST_0),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.h2f_WDATA_0(h2f_WDATA_0),
	.h2f_WDATA_1(h2f_WDATA_1),
	.h2f_WDATA_2(h2f_WDATA_2),
	.h2f_WDATA_3(h2f_WDATA_3),
	.h2f_WDATA_4(h2f_WDATA_4),
	.h2f_WDATA_5(h2f_WDATA_5),
	.h2f_WDATA_6(h2f_WDATA_6),
	.h2f_WDATA_7(h2f_WDATA_7),
	.h2f_WDATA_8(h2f_WDATA_8),
	.h2f_WDATA_9(h2f_WDATA_9),
	.h2f_WDATA_10(h2f_WDATA_10),
	.h2f_WDATA_11(h2f_WDATA_11),
	.h2f_WDATA_12(h2f_WDATA_12),
	.h2f_WDATA_13(h2f_WDATA_13),
	.h2f_WDATA_14(h2f_WDATA_14),
	.h2f_WDATA_15(h2f_WDATA_15),
	.h2f_WDATA_16(h2f_WDATA_16),
	.h2f_WDATA_17(h2f_WDATA_17),
	.h2f_WDATA_18(h2f_WDATA_18),
	.h2f_WDATA_19(h2f_WDATA_19),
	.h2f_WDATA_20(h2f_WDATA_20),
	.h2f_WDATA_21(h2f_WDATA_21),
	.h2f_WDATA_22(h2f_WDATA_22),
	.h2f_WDATA_23(h2f_WDATA_23),
	.h2f_WDATA_24(h2f_WDATA_24),
	.h2f_WDATA_25(h2f_WDATA_25),
	.h2f_WDATA_26(h2f_WDATA_26),
	.h2f_WDATA_27(h2f_WDATA_27),
	.h2f_WDATA_28(h2f_WDATA_28),
	.h2f_WDATA_29(h2f_WDATA_29),
	.h2f_WDATA_30(h2f_WDATA_30),
	.h2f_WDATA_31(h2f_WDATA_31),
	.h2f_WDATA_32(h2f_WDATA_32),
	.h2f_WDATA_33(h2f_WDATA_33),
	.h2f_WDATA_34(h2f_WDATA_34),
	.h2f_WDATA_35(h2f_WDATA_35),
	.h2f_WDATA_36(h2f_WDATA_36),
	.h2f_WDATA_37(h2f_WDATA_37),
	.h2f_WDATA_38(h2f_WDATA_38),
	.h2f_WDATA_39(h2f_WDATA_39),
	.h2f_WDATA_40(h2f_WDATA_40),
	.h2f_WDATA_41(h2f_WDATA_41),
	.h2f_WDATA_42(h2f_WDATA_42),
	.h2f_WDATA_43(h2f_WDATA_43),
	.h2f_WDATA_44(h2f_WDATA_44),
	.h2f_WDATA_45(h2f_WDATA_45),
	.h2f_WDATA_46(h2f_WDATA_46),
	.h2f_WDATA_47(h2f_WDATA_47),
	.h2f_WDATA_48(h2f_WDATA_48),
	.h2f_WDATA_49(h2f_WDATA_49),
	.h2f_WDATA_50(h2f_WDATA_50),
	.h2f_WDATA_51(h2f_WDATA_51),
	.h2f_WDATA_52(h2f_WDATA_52),
	.h2f_WDATA_53(h2f_WDATA_53),
	.h2f_WDATA_54(h2f_WDATA_54),
	.h2f_WDATA_55(h2f_WDATA_55),
	.h2f_WDATA_56(h2f_WDATA_56),
	.h2f_WDATA_57(h2f_WDATA_57),
	.h2f_WDATA_58(h2f_WDATA_58),
	.h2f_WDATA_59(h2f_WDATA_59),
	.h2f_WDATA_60(h2f_WDATA_60),
	.h2f_WDATA_61(h2f_WDATA_61),
	.h2f_WDATA_62(h2f_WDATA_62),
	.h2f_WDATA_63(h2f_WDATA_63),
	.h2f_WDATA_64(h2f_WDATA_64),
	.h2f_WDATA_65(h2f_WDATA_65),
	.h2f_WDATA_66(h2f_WDATA_66),
	.h2f_WDATA_67(h2f_WDATA_67),
	.h2f_WDATA_68(h2f_WDATA_68),
	.h2f_WDATA_69(h2f_WDATA_69),
	.h2f_WDATA_70(h2f_WDATA_70),
	.h2f_WDATA_71(h2f_WDATA_71),
	.h2f_WDATA_72(h2f_WDATA_72),
	.h2f_WDATA_73(h2f_WDATA_73),
	.h2f_WDATA_74(h2f_WDATA_74),
	.h2f_WDATA_75(h2f_WDATA_75),
	.h2f_WDATA_76(h2f_WDATA_76),
	.h2f_WDATA_77(h2f_WDATA_77),
	.h2f_WDATA_78(h2f_WDATA_78),
	.h2f_WDATA_79(h2f_WDATA_79),
	.h2f_WDATA_80(h2f_WDATA_80),
	.h2f_WDATA_81(h2f_WDATA_81),
	.h2f_WDATA_82(h2f_WDATA_82),
	.h2f_WDATA_83(h2f_WDATA_83),
	.h2f_WDATA_84(h2f_WDATA_84),
	.h2f_WDATA_85(h2f_WDATA_85),
	.h2f_WDATA_86(h2f_WDATA_86),
	.h2f_WDATA_87(h2f_WDATA_87),
	.h2f_WDATA_88(h2f_WDATA_88),
	.h2f_WDATA_89(h2f_WDATA_89),
	.h2f_WDATA_90(h2f_WDATA_90),
	.h2f_WDATA_91(h2f_WDATA_91),
	.h2f_WDATA_92(h2f_WDATA_92),
	.h2f_WDATA_93(h2f_WDATA_93),
	.h2f_WDATA_94(h2f_WDATA_94),
	.h2f_WDATA_95(h2f_WDATA_95),
	.h2f_WDATA_96(h2f_WDATA_96),
	.h2f_WDATA_97(h2f_WDATA_97),
	.h2f_WDATA_98(h2f_WDATA_98),
	.h2f_WDATA_99(h2f_WDATA_99),
	.h2f_WDATA_100(h2f_WDATA_100),
	.h2f_WDATA_101(h2f_WDATA_101),
	.h2f_WDATA_102(h2f_WDATA_102),
	.h2f_WDATA_103(h2f_WDATA_103),
	.h2f_WDATA_104(h2f_WDATA_104),
	.h2f_WDATA_105(h2f_WDATA_105),
	.h2f_WDATA_106(h2f_WDATA_106),
	.h2f_WDATA_107(h2f_WDATA_107),
	.h2f_WDATA_108(h2f_WDATA_108),
	.h2f_WDATA_109(h2f_WDATA_109),
	.h2f_WDATA_110(h2f_WDATA_110),
	.h2f_WDATA_111(h2f_WDATA_111),
	.h2f_WDATA_112(h2f_WDATA_112),
	.h2f_WDATA_113(h2f_WDATA_113),
	.h2f_WDATA_114(h2f_WDATA_114),
	.h2f_WDATA_115(h2f_WDATA_115),
	.h2f_WDATA_116(h2f_WDATA_116),
	.h2f_WDATA_117(h2f_WDATA_117),
	.h2f_WDATA_118(h2f_WDATA_118),
	.h2f_WDATA_119(h2f_WDATA_119),
	.h2f_WDATA_120(h2f_WDATA_120),
	.h2f_WDATA_121(h2f_WDATA_121),
	.h2f_WDATA_122(h2f_WDATA_122),
	.h2f_WDATA_123(h2f_WDATA_123),
	.h2f_WDATA_124(h2f_WDATA_124),
	.h2f_WDATA_125(h2f_WDATA_125),
	.h2f_WDATA_126(h2f_WDATA_126),
	.h2f_WDATA_127(h2f_WDATA_127),
	.h2f_WSTRB_0(h2f_WSTRB_0),
	.h2f_WSTRB_1(h2f_WSTRB_1),
	.h2f_WSTRB_2(h2f_WSTRB_2),
	.h2f_WSTRB_3(h2f_WSTRB_3),
	.h2f_WSTRB_4(h2f_WSTRB_4),
	.h2f_WSTRB_5(h2f_WSTRB_5),
	.h2f_WSTRB_6(h2f_WSTRB_6),
	.h2f_WSTRB_7(h2f_WSTRB_7),
	.h2f_WSTRB_8(h2f_WSTRB_8),
	.h2f_WSTRB_9(h2f_WSTRB_9),
	.h2f_WSTRB_10(h2f_WSTRB_10),
	.h2f_WSTRB_11(h2f_WSTRB_11),
	.h2f_WSTRB_12(h2f_WSTRB_12),
	.h2f_WSTRB_13(h2f_WSTRB_13),
	.h2f_WSTRB_14(h2f_WSTRB_14),
	.h2f_WSTRB_15(h2f_WSTRB_15),
	.outclk_wire_0(outclk_wire_0),
	.out_data_37(\fifo_hps_to_fpga_in_cmd_width_adapter|out_data[37]~3_combout ),
	.Mux4(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux4~0_combout ),
	.Mux5(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux5~0_combout ),
	.Mux6(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux6~0_combout ),
	.Mux7(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux7~0_combout ),
	.Mux8(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux8~0_combout ),
	.Mux9(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux9~0_combout ),
	.Mux10(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux10~0_combout ),
	.Mux11(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux11~0_combout ),
	.Mux12(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux12~0_combout ),
	.Mux13(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux13~0_combout ),
	.Mux14(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux14~0_combout ),
	.Mux15(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux15~0_combout ),
	.Mux16(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux16~0_combout ),
	.Mux17(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux17~0_combout ),
	.Mux18(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux18~0_combout ),
	.Mux19(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux19~0_combout ),
	.Mux20(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux20~0_combout ),
	.Mux21(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux21~0_combout ),
	.Mux22(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux22~0_combout ),
	.Mux23(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux23~0_combout ),
	.Mux24(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux24~0_combout ),
	.Mux25(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux25~0_combout ),
	.Mux26(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux26~0_combout ),
	.Mux27(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux27~0_combout ),
	.Mux28(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux28~0_combout ),
	.Mux29(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux29~0_combout ),
	.Mux30(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux30~0_combout ),
	.Mux31(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux31~0_combout ),
	.Mux32(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux32~0_combout ),
	.Mux33(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux33~0_combout ),
	.Mux34(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux34~0_combout ),
	.Mux35(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux35~0_combout ),
	.Mux3(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux3~0_combout ),
	.Mux2(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux2~0_combout ),
	.Mux1(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux1~0_combout ),
	.Mux0(\fifo_hps_to_fpga_in_cmd_width_adapter|Mux0~0_combout ),
	.in_ready_hold(in_ready_hold),
	.Equal0(\router|Equal0~6_combout ),
	.Equal01(\router|Equal0~7_combout ),
	.Equal02(\router|Equal0~14_combout ),
	.nxt_in_ready(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.out_valid_reg(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.count_1(\fifo_hps_to_fpga_in_cmd_width_adapter|count[1]~q ),
	.count_0(\fifo_hps_to_fpga_in_cmd_width_adapter|count[0]~q ),
	.r_sync_rst(r_sync_rst),
	.out_data_2(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[2]~0_combout ),
	.out_data_3(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[3]~1_combout ),
	.src0_valid(\cmd_demux|src0_valid~0_combout ),
	.LessThan2(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|LessThan2~0_combout ),
	.int_output_sel_0(\fifo_hps_to_fpga_in_cmd_width_adapter|int_output_sel[0]~0_combout ),
	.int_output_sel_1(\fifo_hps_to_fpga_in_cmd_width_adapter|int_output_sel[1]~1_combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.src_payload1(\cmd_mux|src_payload~1_combout ),
	.src_payload2(\cmd_mux|src_payload~2_combout ),
	.cp_ready(\fifo_hps_to_fpga_in_agent|cp_ready~1_combout ),
	.out_data_1(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[1]~26_combout ),
	.Decoder0(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|Decoder0~1_combout ),
	.out_data_0(\arm_a9_hps_h2f_axi_master_agent|align_address_to_size|out_data[0]~27_combout ),
	.out_endofpacket(\fifo_hps_to_fpga_in_cmd_width_adapter|out_endofpacket~1_combout ),
	.nxt_in_ready1(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready2(\fifo_hps_to_fpga_in_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.src0_valid1(\cmd_demux|src0_valid~1_combout ),
	.out_data_90(\fifo_hps_to_fpga_in_cmd_width_adapter|out_data[90]~0_combout ),
	.out_data_91(\fifo_hps_to_fpga_in_cmd_width_adapter|out_data[91]~1_combout ),
	.out_data_36(\fifo_hps_to_fpga_in_cmd_width_adapter|out_data[36]~2_combout ));

Computer_System_altera_merlin_width_adapter_3 onchip_sram_s2_rsp_width_adapter(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.q_b_0(q_b_0),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_5(q_b_5),
	.q_b_7(q_b_7),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_21(q_b_21),
	.q_b_23(q_b_23),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.outclk_wire_0(outclk_wire_0),
	.data_reg_0(\onchip_sram_s2_rsp_width_adapter|data_reg[0]~q ),
	.data_reg_1(\onchip_sram_s2_rsp_width_adapter|data_reg[1]~q ),
	.data_reg_2(\onchip_sram_s2_rsp_width_adapter|data_reg[2]~q ),
	.data_reg_3(\onchip_sram_s2_rsp_width_adapter|data_reg[3]~q ),
	.data_reg_4(\onchip_sram_s2_rsp_width_adapter|data_reg[4]~q ),
	.data_reg_5(\onchip_sram_s2_rsp_width_adapter|data_reg[5]~q ),
	.data_reg_6(\onchip_sram_s2_rsp_width_adapter|data_reg[6]~q ),
	.data_reg_7(\onchip_sram_s2_rsp_width_adapter|data_reg[7]~q ),
	.data_reg_8(\onchip_sram_s2_rsp_width_adapter|data_reg[8]~q ),
	.data_reg_9(\onchip_sram_s2_rsp_width_adapter|data_reg[9]~q ),
	.data_reg_10(\onchip_sram_s2_rsp_width_adapter|data_reg[10]~q ),
	.data_reg_11(\onchip_sram_s2_rsp_width_adapter|data_reg[11]~q ),
	.data_reg_12(\onchip_sram_s2_rsp_width_adapter|data_reg[12]~q ),
	.data_reg_13(\onchip_sram_s2_rsp_width_adapter|data_reg[13]~q ),
	.data_reg_14(\onchip_sram_s2_rsp_width_adapter|data_reg[14]~q ),
	.data_reg_15(\onchip_sram_s2_rsp_width_adapter|data_reg[15]~q ),
	.data_reg_16(\onchip_sram_s2_rsp_width_adapter|data_reg[16]~q ),
	.data_reg_17(\onchip_sram_s2_rsp_width_adapter|data_reg[17]~q ),
	.data_reg_18(\onchip_sram_s2_rsp_width_adapter|data_reg[18]~q ),
	.data_reg_19(\onchip_sram_s2_rsp_width_adapter|data_reg[19]~q ),
	.data_reg_20(\onchip_sram_s2_rsp_width_adapter|data_reg[20]~q ),
	.data_reg_21(\onchip_sram_s2_rsp_width_adapter|data_reg[21]~q ),
	.data_reg_22(\onchip_sram_s2_rsp_width_adapter|data_reg[22]~q ),
	.data_reg_23(\onchip_sram_s2_rsp_width_adapter|data_reg[23]~q ),
	.data_reg_24(\onchip_sram_s2_rsp_width_adapter|data_reg[24]~q ),
	.data_reg_25(\onchip_sram_s2_rsp_width_adapter|data_reg[25]~q ),
	.data_reg_26(\onchip_sram_s2_rsp_width_adapter|data_reg[26]~q ),
	.data_reg_27(\onchip_sram_s2_rsp_width_adapter|data_reg[27]~q ),
	.data_reg_28(\onchip_sram_s2_rsp_width_adapter|data_reg[28]~q ),
	.data_reg_29(\onchip_sram_s2_rsp_width_adapter|data_reg[29]~q ),
	.data_reg_30(\onchip_sram_s2_rsp_width_adapter|data_reg[30]~q ),
	.data_reg_31(\onchip_sram_s2_rsp_width_adapter|data_reg[31]~q ),
	.data_reg_32(\onchip_sram_s2_rsp_width_adapter|data_reg[32]~q ),
	.data_reg_33(\onchip_sram_s2_rsp_width_adapter|data_reg[33]~q ),
	.data_reg_34(\onchip_sram_s2_rsp_width_adapter|data_reg[34]~q ),
	.data_reg_35(\onchip_sram_s2_rsp_width_adapter|data_reg[35]~q ),
	.data_reg_36(\onchip_sram_s2_rsp_width_adapter|data_reg[36]~q ),
	.data_reg_37(\onchip_sram_s2_rsp_width_adapter|data_reg[37]~q ),
	.data_reg_38(\onchip_sram_s2_rsp_width_adapter|data_reg[38]~q ),
	.data_reg_39(\onchip_sram_s2_rsp_width_adapter|data_reg[39]~q ),
	.data_reg_40(\onchip_sram_s2_rsp_width_adapter|data_reg[40]~q ),
	.data_reg_41(\onchip_sram_s2_rsp_width_adapter|data_reg[41]~q ),
	.data_reg_42(\onchip_sram_s2_rsp_width_adapter|data_reg[42]~q ),
	.data_reg_43(\onchip_sram_s2_rsp_width_adapter|data_reg[43]~q ),
	.data_reg_44(\onchip_sram_s2_rsp_width_adapter|data_reg[44]~q ),
	.data_reg_45(\onchip_sram_s2_rsp_width_adapter|data_reg[45]~q ),
	.data_reg_46(\onchip_sram_s2_rsp_width_adapter|data_reg[46]~q ),
	.data_reg_47(\onchip_sram_s2_rsp_width_adapter|data_reg[47]~q ),
	.data_reg_48(\onchip_sram_s2_rsp_width_adapter|data_reg[48]~q ),
	.data_reg_49(\onchip_sram_s2_rsp_width_adapter|data_reg[49]~q ),
	.data_reg_50(\onchip_sram_s2_rsp_width_adapter|data_reg[50]~q ),
	.data_reg_51(\onchip_sram_s2_rsp_width_adapter|data_reg[51]~q ),
	.data_reg_52(\onchip_sram_s2_rsp_width_adapter|data_reg[52]~q ),
	.data_reg_53(\onchip_sram_s2_rsp_width_adapter|data_reg[53]~q ),
	.data_reg_54(\onchip_sram_s2_rsp_width_adapter|data_reg[54]~q ),
	.data_reg_55(\onchip_sram_s2_rsp_width_adapter|data_reg[55]~q ),
	.data_reg_56(\onchip_sram_s2_rsp_width_adapter|data_reg[56]~q ),
	.data_reg_57(\onchip_sram_s2_rsp_width_adapter|data_reg[57]~q ),
	.data_reg_58(\onchip_sram_s2_rsp_width_adapter|data_reg[58]~q ),
	.data_reg_59(\onchip_sram_s2_rsp_width_adapter|data_reg[59]~q ),
	.data_reg_60(\onchip_sram_s2_rsp_width_adapter|data_reg[60]~q ),
	.data_reg_61(\onchip_sram_s2_rsp_width_adapter|data_reg[61]~q ),
	.data_reg_62(\onchip_sram_s2_rsp_width_adapter|data_reg[62]~q ),
	.data_reg_63(\onchip_sram_s2_rsp_width_adapter|data_reg[63]~q ),
	.data_reg_64(\onchip_sram_s2_rsp_width_adapter|data_reg[64]~q ),
	.data_reg_65(\onchip_sram_s2_rsp_width_adapter|data_reg[65]~q ),
	.data_reg_66(\onchip_sram_s2_rsp_width_adapter|data_reg[66]~q ),
	.data_reg_67(\onchip_sram_s2_rsp_width_adapter|data_reg[67]~q ),
	.data_reg_68(\onchip_sram_s2_rsp_width_adapter|data_reg[68]~q ),
	.data_reg_69(\onchip_sram_s2_rsp_width_adapter|data_reg[69]~q ),
	.data_reg_70(\onchip_sram_s2_rsp_width_adapter|data_reg[70]~q ),
	.data_reg_71(\onchip_sram_s2_rsp_width_adapter|data_reg[71]~q ),
	.data_reg_72(\onchip_sram_s2_rsp_width_adapter|data_reg[72]~q ),
	.data_reg_73(\onchip_sram_s2_rsp_width_adapter|data_reg[73]~q ),
	.data_reg_74(\onchip_sram_s2_rsp_width_adapter|data_reg[74]~q ),
	.data_reg_75(\onchip_sram_s2_rsp_width_adapter|data_reg[75]~q ),
	.data_reg_76(\onchip_sram_s2_rsp_width_adapter|data_reg[76]~q ),
	.data_reg_77(\onchip_sram_s2_rsp_width_adapter|data_reg[77]~q ),
	.data_reg_78(\onchip_sram_s2_rsp_width_adapter|data_reg[78]~q ),
	.data_reg_79(\onchip_sram_s2_rsp_width_adapter|data_reg[79]~q ),
	.data_reg_80(\onchip_sram_s2_rsp_width_adapter|data_reg[80]~q ),
	.data_reg_81(\onchip_sram_s2_rsp_width_adapter|data_reg[81]~q ),
	.data_reg_82(\onchip_sram_s2_rsp_width_adapter|data_reg[82]~q ),
	.data_reg_83(\onchip_sram_s2_rsp_width_adapter|data_reg[83]~q ),
	.data_reg_84(\onchip_sram_s2_rsp_width_adapter|data_reg[84]~q ),
	.data_reg_85(\onchip_sram_s2_rsp_width_adapter|data_reg[85]~q ),
	.data_reg_86(\onchip_sram_s2_rsp_width_adapter|data_reg[86]~q ),
	.data_reg_87(\onchip_sram_s2_rsp_width_adapter|data_reg[87]~q ),
	.data_reg_88(\onchip_sram_s2_rsp_width_adapter|data_reg[88]~q ),
	.data_reg_89(\onchip_sram_s2_rsp_width_adapter|data_reg[89]~q ),
	.data_reg_90(\onchip_sram_s2_rsp_width_adapter|data_reg[90]~q ),
	.data_reg_91(\onchip_sram_s2_rsp_width_adapter|data_reg[91]~q ),
	.data_reg_92(\onchip_sram_s2_rsp_width_adapter|data_reg[92]~q ),
	.data_reg_93(\onchip_sram_s2_rsp_width_adapter|data_reg[93]~q ),
	.data_reg_94(\onchip_sram_s2_rsp_width_adapter|data_reg[94]~q ),
	.data_reg_95(\onchip_sram_s2_rsp_width_adapter|data_reg[95]~q ),
	.read_latency_shift_reg_0(\onchip_sram_s2_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\onchip_sram_s2_agent_rdata_fifo|mem_used[0]~q ),
	.mem_125_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][125]~q ),
	.mem_used_01(\onchip_sram_s2_agent_rsp_fifo|mem_used[0]~q ),
	.out_valid(\onchip_sram_s2_rsp_width_adapter|out_valid~0_combout ),
	.comb(\onchip_sram_s2_agent|comb~0_combout ),
	.burst_uncompress_busy(\onchip_sram_s2_agent|uncompressor|burst_uncompress_busy~q ),
	.src_payload(\rsp_mux_001|src_payload~0_combout ),
	.mem_38_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][38]~q ),
	.source_addr_2(\onchip_sram_s2_agent|uncompressor|source_addr[2]~0_combout ),
	.source_addr_21(\onchip_sram_s2_agent|uncompressor|source_addr[2]~1_combout ),
	.mem_122_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][122]~q ),
	.mem_123_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][123]~q ),
	.mem_91_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][91]~q ),
	.mem_124_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][124]~q ),
	.mem_90_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][90]~q ),
	.mem_39_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][39]~q ),
	.source_addr_3(\onchip_sram_s2_agent|uncompressor|source_addr[3]~2_combout ),
	.always10(\onchip_sram_s2_rsp_width_adapter|always10~9_combout ),
	.src0_valid(\rsp_demux_001|src0_valid~0_combout ),
	.ShiftLeft0(\onchip_sram_s2_rsp_width_adapter|ShiftLeft0~0_combout ),
	.always4(\onchip_sram_s2_agent_rdata_fifo|always4~0_combout ),
	.mem_0_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][0]~q ),
	.LessThan15(\onchip_sram_s2_rsp_width_adapter|LessThan15~0_combout ),
	.mem_2_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][2]~q ),
	.mem_3_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][3]~q ),
	.mem_5_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][5]~q ),
	.mem_7_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][7]~q ),
	.mem_9_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][9]~q ),
	.mem_10_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][10]~q ),
	.mem_11_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][11]~q ),
	.mem_12_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][12]~q ),
	.mem_14_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][14]~q ),
	.mem_15_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][15]~q ),
	.mem_16_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][16]~q ),
	.mem_18_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][18]~q ),
	.mem_19_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][19]~q ),
	.mem_21_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][21]~q ),
	.mem_23_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][23]~q ),
	.mem_25_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][25]~q ),
	.mem_26_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][26]~q ),
	.mem_27_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][27]~q ),
	.mem_28_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][28]~q ),
	.mem_30_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][30]~q ),
	.mem_31_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][31]~q ),
	.ShiftLeft01(\onchip_sram_s2_rsp_width_adapter|ShiftLeft0~1_combout ),
	.ShiftLeft02(\onchip_sram_s2_rsp_width_adapter|ShiftLeft0~2_combout ),
	.out_data_1(\onchip_sram_s2_agent_rdata_fifo|out_data[1]~0_combout ),
	.out_data_4(\onchip_sram_s2_agent_rdata_fifo|out_data[4]~1_combout ),
	.out_data_6(\onchip_sram_s2_agent_rdata_fifo|out_data[6]~2_combout ),
	.out_data_8(\onchip_sram_s2_agent_rdata_fifo|out_data[8]~3_combout ),
	.out_data_13(\onchip_sram_s2_agent_rdata_fifo|out_data[13]~4_combout ),
	.out_data_17(\onchip_sram_s2_agent_rdata_fifo|out_data[17]~5_combout ),
	.out_data_20(\onchip_sram_s2_agent_rdata_fifo|out_data[20]~6_combout ),
	.out_data_22(\onchip_sram_s2_agent_rdata_fifo|out_data[22]~7_combout ),
	.out_data_24(\onchip_sram_s2_agent_rdata_fifo|out_data[24]~8_combout ),
	.out_data_29(\onchip_sram_s2_agent_rdata_fifo|out_data[29]~9_combout ),
	.r_sync_rst(r_sync_rst),
	.p1_ready(\onchip_sram_s2_rsp_width_adapter|p1_ready~0_combout ),
	.always101(\onchip_sram_s2_rsp_width_adapter|always10~10_combout ));

Computer_System_altera_merlin_width_adapter_1 fifo_hps_to_fpga_in_rsp_width_adapter(
	.h2f_BREADY_0(h2f_BREADY_0),
	.h2f_RREADY_0(h2f_RREADY_0),
	.outclk_wire_0(outclk_wire_0),
	.data_reg_0(\fifo_hps_to_fpga_in_rsp_width_adapter|data_reg[0]~q ),
	.data_reg_32(\fifo_hps_to_fpga_in_rsp_width_adapter|data_reg[32]~q ),
	.data_reg_64(\fifo_hps_to_fpga_in_rsp_width_adapter|data_reg[64]~q ),
	.mem_68_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][68]~q ),
	.mem_122_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][122]~q ),
	.mem_123_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][123]~q ),
	.mem_124_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][124]~q ),
	.mem_90_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][90]~q ),
	.mem_91_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][91]~q ),
	.ShiftRight0(\fifo_hps_to_fpga_in_rsp_width_adapter|ShiftRight0~0_combout ),
	.source_addr_2(\fifo_hps_to_fpga_in_agent|uncompressor|source_addr[2]~0_combout ),
	.always10(\fifo_hps_to_fpga_in_rsp_width_adapter|always10~0_combout ),
	.mem_126_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][126]~q ),
	.source_addr_3(\fifo_hps_to_fpga_in_agent|uncompressor|source_addr[3]~1_combout ),
	.always101(\fifo_hps_to_fpga_in_rsp_width_adapter|always10~1_combout ),
	.mem_31_0(\fifo_hps_to_fpga_in_agent_rdata_fifo|mem[0][31]~q ),
	.LessThan15(\fifo_hps_to_fpga_in_rsp_width_adapter|LessThan15~0_combout ),
	.r_sync_rst(r_sync_rst),
	.p1_ready(\fifo_hps_to_fpga_in_rsp_width_adapter|p1_ready~0_combout ),
	.read(\fifo_hps_to_fpga_in_agent_rsp_fifo|read~0_combout ),
	.always102(\fifo_hps_to_fpga_in_rsp_width_adapter|always10~2_combout ));

Computer_System_Computer_System_mm_interconnect_0_rsp_mux_1 rsp_mux_001(
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.data_reg_0(\fifo_hps_to_fpga_in_rsp_width_adapter|data_reg[0]~q ),
	.data_reg_01(\onchip_sram_s2_rsp_width_adapter|data_reg[0]~q ),
	.data_reg_1(\onchip_sram_s2_rsp_width_adapter|data_reg[1]~q ),
	.data_reg_2(\onchip_sram_s2_rsp_width_adapter|data_reg[2]~q ),
	.data_reg_3(\onchip_sram_s2_rsp_width_adapter|data_reg[3]~q ),
	.data_reg_4(\onchip_sram_s2_rsp_width_adapter|data_reg[4]~q ),
	.data_reg_5(\onchip_sram_s2_rsp_width_adapter|data_reg[5]~q ),
	.data_reg_6(\onchip_sram_s2_rsp_width_adapter|data_reg[6]~q ),
	.data_reg_7(\onchip_sram_s2_rsp_width_adapter|data_reg[7]~q ),
	.data_reg_8(\onchip_sram_s2_rsp_width_adapter|data_reg[8]~q ),
	.data_reg_9(\onchip_sram_s2_rsp_width_adapter|data_reg[9]~q ),
	.data_reg_10(\onchip_sram_s2_rsp_width_adapter|data_reg[10]~q ),
	.data_reg_11(\onchip_sram_s2_rsp_width_adapter|data_reg[11]~q ),
	.data_reg_12(\onchip_sram_s2_rsp_width_adapter|data_reg[12]~q ),
	.data_reg_13(\onchip_sram_s2_rsp_width_adapter|data_reg[13]~q ),
	.data_reg_14(\onchip_sram_s2_rsp_width_adapter|data_reg[14]~q ),
	.data_reg_15(\onchip_sram_s2_rsp_width_adapter|data_reg[15]~q ),
	.data_reg_16(\onchip_sram_s2_rsp_width_adapter|data_reg[16]~q ),
	.data_reg_17(\onchip_sram_s2_rsp_width_adapter|data_reg[17]~q ),
	.data_reg_18(\onchip_sram_s2_rsp_width_adapter|data_reg[18]~q ),
	.data_reg_19(\onchip_sram_s2_rsp_width_adapter|data_reg[19]~q ),
	.data_reg_20(\onchip_sram_s2_rsp_width_adapter|data_reg[20]~q ),
	.data_reg_21(\onchip_sram_s2_rsp_width_adapter|data_reg[21]~q ),
	.data_reg_22(\onchip_sram_s2_rsp_width_adapter|data_reg[22]~q ),
	.data_reg_23(\onchip_sram_s2_rsp_width_adapter|data_reg[23]~q ),
	.data_reg_24(\onchip_sram_s2_rsp_width_adapter|data_reg[24]~q ),
	.data_reg_25(\onchip_sram_s2_rsp_width_adapter|data_reg[25]~q ),
	.data_reg_26(\onchip_sram_s2_rsp_width_adapter|data_reg[26]~q ),
	.data_reg_27(\onchip_sram_s2_rsp_width_adapter|data_reg[27]~q ),
	.data_reg_28(\onchip_sram_s2_rsp_width_adapter|data_reg[28]~q ),
	.data_reg_29(\onchip_sram_s2_rsp_width_adapter|data_reg[29]~q ),
	.data_reg_30(\onchip_sram_s2_rsp_width_adapter|data_reg[30]~q ),
	.data_reg_31(\onchip_sram_s2_rsp_width_adapter|data_reg[31]~q ),
	.data_reg_32(\fifo_hps_to_fpga_in_rsp_width_adapter|data_reg[32]~q ),
	.data_reg_321(\onchip_sram_s2_rsp_width_adapter|data_reg[32]~q ),
	.data_reg_33(\onchip_sram_s2_rsp_width_adapter|data_reg[33]~q ),
	.data_reg_34(\onchip_sram_s2_rsp_width_adapter|data_reg[34]~q ),
	.data_reg_35(\onchip_sram_s2_rsp_width_adapter|data_reg[35]~q ),
	.data_reg_36(\onchip_sram_s2_rsp_width_adapter|data_reg[36]~q ),
	.data_reg_37(\onchip_sram_s2_rsp_width_adapter|data_reg[37]~q ),
	.data_reg_38(\onchip_sram_s2_rsp_width_adapter|data_reg[38]~q ),
	.data_reg_39(\onchip_sram_s2_rsp_width_adapter|data_reg[39]~q ),
	.data_reg_40(\onchip_sram_s2_rsp_width_adapter|data_reg[40]~q ),
	.data_reg_41(\onchip_sram_s2_rsp_width_adapter|data_reg[41]~q ),
	.data_reg_42(\onchip_sram_s2_rsp_width_adapter|data_reg[42]~q ),
	.data_reg_43(\onchip_sram_s2_rsp_width_adapter|data_reg[43]~q ),
	.data_reg_44(\onchip_sram_s2_rsp_width_adapter|data_reg[44]~q ),
	.data_reg_45(\onchip_sram_s2_rsp_width_adapter|data_reg[45]~q ),
	.data_reg_46(\onchip_sram_s2_rsp_width_adapter|data_reg[46]~q ),
	.data_reg_47(\onchip_sram_s2_rsp_width_adapter|data_reg[47]~q ),
	.data_reg_48(\onchip_sram_s2_rsp_width_adapter|data_reg[48]~q ),
	.data_reg_49(\onchip_sram_s2_rsp_width_adapter|data_reg[49]~q ),
	.data_reg_50(\onchip_sram_s2_rsp_width_adapter|data_reg[50]~q ),
	.data_reg_51(\onchip_sram_s2_rsp_width_adapter|data_reg[51]~q ),
	.data_reg_52(\onchip_sram_s2_rsp_width_adapter|data_reg[52]~q ),
	.data_reg_53(\onchip_sram_s2_rsp_width_adapter|data_reg[53]~q ),
	.data_reg_54(\onchip_sram_s2_rsp_width_adapter|data_reg[54]~q ),
	.data_reg_55(\onchip_sram_s2_rsp_width_adapter|data_reg[55]~q ),
	.data_reg_56(\onchip_sram_s2_rsp_width_adapter|data_reg[56]~q ),
	.data_reg_57(\onchip_sram_s2_rsp_width_adapter|data_reg[57]~q ),
	.data_reg_58(\onchip_sram_s2_rsp_width_adapter|data_reg[58]~q ),
	.data_reg_59(\onchip_sram_s2_rsp_width_adapter|data_reg[59]~q ),
	.data_reg_60(\onchip_sram_s2_rsp_width_adapter|data_reg[60]~q ),
	.data_reg_61(\onchip_sram_s2_rsp_width_adapter|data_reg[61]~q ),
	.data_reg_62(\onchip_sram_s2_rsp_width_adapter|data_reg[62]~q ),
	.data_reg_63(\onchip_sram_s2_rsp_width_adapter|data_reg[63]~q ),
	.data_reg_64(\fifo_hps_to_fpga_in_rsp_width_adapter|data_reg[64]~q ),
	.data_reg_641(\onchip_sram_s2_rsp_width_adapter|data_reg[64]~q ),
	.data_reg_65(\onchip_sram_s2_rsp_width_adapter|data_reg[65]~q ),
	.data_reg_66(\onchip_sram_s2_rsp_width_adapter|data_reg[66]~q ),
	.data_reg_67(\onchip_sram_s2_rsp_width_adapter|data_reg[67]~q ),
	.data_reg_68(\onchip_sram_s2_rsp_width_adapter|data_reg[68]~q ),
	.data_reg_69(\onchip_sram_s2_rsp_width_adapter|data_reg[69]~q ),
	.data_reg_70(\onchip_sram_s2_rsp_width_adapter|data_reg[70]~q ),
	.data_reg_71(\onchip_sram_s2_rsp_width_adapter|data_reg[71]~q ),
	.data_reg_72(\onchip_sram_s2_rsp_width_adapter|data_reg[72]~q ),
	.data_reg_73(\onchip_sram_s2_rsp_width_adapter|data_reg[73]~q ),
	.data_reg_74(\onchip_sram_s2_rsp_width_adapter|data_reg[74]~q ),
	.data_reg_75(\onchip_sram_s2_rsp_width_adapter|data_reg[75]~q ),
	.data_reg_76(\onchip_sram_s2_rsp_width_adapter|data_reg[76]~q ),
	.data_reg_77(\onchip_sram_s2_rsp_width_adapter|data_reg[77]~q ),
	.data_reg_78(\onchip_sram_s2_rsp_width_adapter|data_reg[78]~q ),
	.data_reg_79(\onchip_sram_s2_rsp_width_adapter|data_reg[79]~q ),
	.data_reg_80(\onchip_sram_s2_rsp_width_adapter|data_reg[80]~q ),
	.data_reg_81(\onchip_sram_s2_rsp_width_adapter|data_reg[81]~q ),
	.data_reg_82(\onchip_sram_s2_rsp_width_adapter|data_reg[82]~q ),
	.data_reg_83(\onchip_sram_s2_rsp_width_adapter|data_reg[83]~q ),
	.data_reg_84(\onchip_sram_s2_rsp_width_adapter|data_reg[84]~q ),
	.data_reg_85(\onchip_sram_s2_rsp_width_adapter|data_reg[85]~q ),
	.data_reg_86(\onchip_sram_s2_rsp_width_adapter|data_reg[86]~q ),
	.data_reg_87(\onchip_sram_s2_rsp_width_adapter|data_reg[87]~q ),
	.data_reg_88(\onchip_sram_s2_rsp_width_adapter|data_reg[88]~q ),
	.data_reg_89(\onchip_sram_s2_rsp_width_adapter|data_reg[89]~q ),
	.data_reg_90(\onchip_sram_s2_rsp_width_adapter|data_reg[90]~q ),
	.data_reg_91(\onchip_sram_s2_rsp_width_adapter|data_reg[91]~q ),
	.data_reg_92(\onchip_sram_s2_rsp_width_adapter|data_reg[92]~q ),
	.data_reg_93(\onchip_sram_s2_rsp_width_adapter|data_reg[93]~q ),
	.data_reg_94(\onchip_sram_s2_rsp_width_adapter|data_reg[94]~q ),
	.data_reg_95(\onchip_sram_s2_rsp_width_adapter|data_reg[95]~q ),
	.out_valid(\onchip_sram_s2_rsp_width_adapter|out_valid~0_combout ),
	.comb(\onchip_sram_s2_agent|comb~0_combout ),
	.mem_126_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][126]~q ),
	.mem_66_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][66]~q ),
	.burst_uncompress_busy(\onchip_sram_s2_agent|uncompressor|burst_uncompress_busy~q ),
	.last_packet_beat(\onchip_sram_s2_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat1(\onchip_sram_s2_agent|uncompressor|last_packet_beat~1_combout ),
	.last_packet_beat2(\onchip_sram_s2_agent|uncompressor|last_packet_beat~4_combout ),
	.src_payload(\rsp_mux_001|src_payload~0_combout ),
	.mem_38_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][38]~q ),
	.source_addr_2(\onchip_sram_s2_agent|uncompressor|source_addr[2]~0_combout ),
	.mem_39_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][39]~q ),
	.source_addr_3(\onchip_sram_s2_agent|uncompressor|source_addr[3]~2_combout ),
	.always10(\onchip_sram_s2_rsp_width_adapter|always10~9_combout ),
	.src0_valid(\rsp_demux_001|src0_valid~0_combout ),
	.mem_68_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][68]~q ),
	.comb1(\fifo_hps_to_fpga_in_agent|comb~0_combout ),
	.ShiftRight0(\fifo_hps_to_fpga_in_rsp_width_adapter|ShiftRight0~0_combout ),
	.source_addr_21(\fifo_hps_to_fpga_in_agent|uncompressor|source_addr[2]~0_combout ),
	.always101(\fifo_hps_to_fpga_in_rsp_width_adapter|always10~0_combout ),
	.mem_126_01(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][126]~q ),
	.source_addr_31(\fifo_hps_to_fpga_in_agent|uncompressor|source_addr[3]~1_combout ),
	.always102(\fifo_hps_to_fpga_in_rsp_width_adapter|always10~1_combout ),
	.src_payload_0(src_payload_0),
	.src1_valid(\rsp_demux|src1_valid~0_combout ),
	.WideOr11(WideOr11),
	.mem_101_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][101]~q ),
	.mem_101_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][101]~q ),
	.mem_102_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][102]~q ),
	.mem_102_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][102]~q ),
	.mem_103_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][103]~q ),
	.mem_103_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][103]~q ),
	.mem_104_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][104]~q ),
	.mem_104_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][104]~q ),
	.mem_105_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][105]~q ),
	.mem_106_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][106]~q ),
	.mem_107_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][107]~q ),
	.mem_108_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][108]~q ),
	.mem_109_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][109]~q ),
	.mem_110_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][110]~q ),
	.mem_111_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][111]~q ),
	.mem_112_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][112]~q ),
	.mem_31_0(\fifo_hps_to_fpga_in_agent_rdata_fifo|mem[0][31]~q ),
	.LessThan15(\fifo_hps_to_fpga_in_rsp_width_adapter|LessThan15~0_combout ),
	.ShiftLeft0(\onchip_sram_s2_rsp_width_adapter|ShiftLeft0~0_combout ),
	.always4(\onchip_sram_s2_agent_rdata_fifo|always4~0_combout ),
	.mem_0_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][0]~q ),
	.LessThan151(\onchip_sram_s2_rsp_width_adapter|LessThan15~0_combout ),
	.src_data_0(src_data_0),
	.mem_1_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][1]~q ),
	.src_payload1(src_payload),
	.mem_2_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][2]~q ),
	.src_data_2(src_data_2),
	.mem_3_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][3]~q ),
	.src_data_3(src_data_3),
	.mem_4_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][4]~q ),
	.src_payload2(src_payload1),
	.mem_5_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][5]~q ),
	.src_data_5(src_data_5),
	.mem_6_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][6]~q ),
	.src_payload3(src_payload2),
	.mem_7_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][7]~q ),
	.src_data_7(src_data_7),
	.mem_8_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][8]~q ),
	.src_payload4(src_payload3),
	.mem_9_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][9]~q ),
	.src_data_9(src_data_9),
	.mem_10_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][10]~q ),
	.src_data_10(src_data_10),
	.mem_11_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][11]~q ),
	.src_data_11(src_data_11),
	.mem_12_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][12]~q ),
	.src_data_12(src_data_12),
	.mem_13_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][13]~q ),
	.src_payload5(src_payload4),
	.mem_14_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][14]~q ),
	.src_data_14(src_data_14),
	.mem_15_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][15]~q ),
	.src_data_15(src_data_15),
	.mem_16_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][16]~q ),
	.src_data_16(src_data_16),
	.mem_17_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][17]~q ),
	.src_payload6(src_payload5),
	.mem_18_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][18]~q ),
	.src_data_18(src_data_18),
	.mem_19_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][19]~q ),
	.src_data_19(src_data_19),
	.mem_20_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][20]~q ),
	.src_payload7(src_payload6),
	.mem_21_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][21]~q ),
	.src_data_21(src_data_21),
	.mem_22_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][22]~q ),
	.src_payload8(src_payload7),
	.mem_23_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][23]~q ),
	.src_data_23(src_data_23),
	.mem_24_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][24]~q ),
	.src_payload9(src_payload8),
	.mem_25_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][25]~q ),
	.src_data_25(src_data_25),
	.mem_26_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][26]~q ),
	.src_data_26(src_data_26),
	.mem_27_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][27]~q ),
	.src_data_27(src_data_27),
	.mem_28_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][28]~q ),
	.src_data_28(src_data_28),
	.mem_29_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][29]~q ),
	.src_payload10(src_payload9),
	.mem_30_0(\onchip_sram_s2_agent_rdata_fifo|mem[0][30]~q ),
	.src_data_30(src_data_30),
	.mem_31_01(\onchip_sram_s2_agent_rdata_fifo|mem[0][31]~q ),
	.src_data_31(src_data_31),
	.ShiftLeft01(\onchip_sram_s2_rsp_width_adapter|ShiftLeft0~1_combout ),
	.src_data_32(src_data_32),
	.src_payload11(src_payload10),
	.src_data_34(src_data_34),
	.src_data_35(src_data_35),
	.src_payload12(src_payload11),
	.src_data_37(src_data_37),
	.src_payload13(src_payload12),
	.src_data_39(src_data_39),
	.src_payload14(src_payload13),
	.src_data_41(src_data_41),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_payload15(src_payload14),
	.src_data_46(src_data_46),
	.src_data_47(src_data_47),
	.src_data_48(src_data_48),
	.src_payload16(src_payload15),
	.src_data_50(src_data_50),
	.src_data_51(src_data_51),
	.src_payload17(src_payload16),
	.src_data_53(src_data_53),
	.src_payload18(src_payload17),
	.src_data_55(src_data_55),
	.src_payload19(src_payload18),
	.src_data_57(src_data_57),
	.src_data_58(src_data_58),
	.src_data_59(src_data_59),
	.src_data_60(src_data_60),
	.src_payload20(src_payload19),
	.src_data_62(src_data_62),
	.src_data_63(src_data_63),
	.ShiftLeft02(\onchip_sram_s2_rsp_width_adapter|ShiftLeft0~2_combout ),
	.src_data_64(src_data_64),
	.src_payload21(src_payload20),
	.src_data_66(src_data_66),
	.src_data_67(src_data_67),
	.src_payload22(src_payload21),
	.src_data_69(src_data_69),
	.src_payload23(src_payload22),
	.src_data_71(src_data_71),
	.src_payload24(src_payload23),
	.src_data_73(src_data_73),
	.src_data_74(src_data_74),
	.src_data_75(src_data_75),
	.src_data_76(src_data_76),
	.src_payload25(src_payload24),
	.src_data_78(src_data_78),
	.src_data_79(src_data_79),
	.src_data_80(src_data_80),
	.src_payload26(src_payload25),
	.src_data_82(src_data_82),
	.src_data_83(src_data_83),
	.src_payload27(src_payload26),
	.src_data_85(src_data_85),
	.src_payload28(src_payload27),
	.src_data_87(src_data_87),
	.src_payload29(src_payload28),
	.src_data_89(src_data_89),
	.src_data_90(src_data_90),
	.src_data_91(src_data_91),
	.src_data_92(src_data_92),
	.src_payload30(src_payload29),
	.src_data_94(src_data_94),
	.src_data_95(src_data_95),
	.src_data_96(src_data_96),
	.out_data_1(\onchip_sram_s2_agent_rdata_fifo|out_data[1]~0_combout ),
	.src_payload31(src_payload30),
	.src_data_98(src_data_98),
	.src_data_99(src_data_99),
	.out_data_4(\onchip_sram_s2_agent_rdata_fifo|out_data[4]~1_combout ),
	.src_payload32(src_payload31),
	.src_data_101(src_data_101),
	.out_data_6(\onchip_sram_s2_agent_rdata_fifo|out_data[6]~2_combout ),
	.src_payload33(src_payload32),
	.src_data_103(src_data_103),
	.out_data_8(\onchip_sram_s2_agent_rdata_fifo|out_data[8]~3_combout ),
	.src_payload34(src_payload33),
	.src_data_105(src_data_105),
	.src_data_106(src_data_106),
	.src_data_107(src_data_107),
	.src_data_108(src_data_108),
	.out_data_13(\onchip_sram_s2_agent_rdata_fifo|out_data[13]~4_combout ),
	.src_payload35(src_payload34),
	.src_data_110(src_data_110),
	.src_data_111(src_data_111),
	.src_data_112(src_data_112),
	.out_data_17(\onchip_sram_s2_agent_rdata_fifo|out_data[17]~5_combout ),
	.src_payload36(src_payload35),
	.src_data_114(src_data_114),
	.src_data_115(src_data_115),
	.out_data_20(\onchip_sram_s2_agent_rdata_fifo|out_data[20]~6_combout ),
	.src_payload37(src_payload36),
	.src_data_117(src_data_117),
	.out_data_22(\onchip_sram_s2_agent_rdata_fifo|out_data[22]~7_combout ),
	.src_payload38(src_payload37),
	.src_data_119(src_data_119),
	.out_data_24(\onchip_sram_s2_agent_rdata_fifo|out_data[24]~8_combout ),
	.src_payload39(src_payload38),
	.src_data_121(src_data_121),
	.src_data_122(src_data_122),
	.src_data_123(src_data_123),
	.src_data_124(src_data_124),
	.out_data_29(\onchip_sram_s2_agent_rdata_fifo|out_data[29]~9_combout ),
	.src_payload40(src_payload39),
	.src_data_126(src_data_126),
	.src_data_127(src_data_127),
	.src_data_209(src_data_2091),
	.src_data_210(src_data_2101),
	.src_data_211(src_data_2111),
	.src_data_212(src_data_2121),
	.src_data_213(src_data_2131),
	.src_data_214(src_data_2141),
	.src_data_215(src_data_2151),
	.src_data_216(src_data_2161),
	.src_data_217(src_data_2171),
	.src_data_218(src_data_2181),
	.src_data_219(src_data_2191),
	.src_data_220(src_data_2201),
	.src_payload41(\rsp_mux_001|src_payload~93_combout ));

Computer_System_Computer_System_mm_interconnect_0_rsp_mux rsp_mux(
	.out_valid(\onchip_sram_s2_rsp_width_adapter|out_valid~0_combout ),
	.src_payload(\rsp_mux_001|src_payload~0_combout ),
	.always10(\onchip_sram_s2_rsp_width_adapter|always10~9_combout ),
	.src0_valid(\rsp_demux_001|src0_valid~0_combout ),
	.mem_68_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][68]~q ),
	.comb(\fifo_hps_to_fpga_in_agent|comb~0_combout ),
	.ShiftRight0(\fifo_hps_to_fpga_in_rsp_width_adapter|ShiftRight0~0_combout ),
	.always101(\fifo_hps_to_fpga_in_rsp_width_adapter|always10~0_combout ),
	.always102(\fifo_hps_to_fpga_in_rsp_width_adapter|always10~1_combout ),
	.src0_valid1(\rsp_demux|src0_valid~0_combout ),
	.WideOr11(WideOr1),
	.mem_101_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][101]~q ),
	.mem_101_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][101]~q ),
	.src_data_209(src_data_209),
	.mem_102_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][102]~q ),
	.mem_102_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][102]~q ),
	.src_data_210(src_data_210),
	.mem_103_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][103]~q ),
	.mem_103_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][103]~q ),
	.src_data_211(src_data_211),
	.mem_104_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][104]~q ),
	.mem_104_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][104]~q ),
	.src_data_212(src_data_212),
	.mem_105_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][105]~q ),
	.mem_105_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][105]~q ),
	.src_data_213(src_data_213),
	.mem_106_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][106]~q ),
	.mem_106_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][106]~q ),
	.src_data_214(src_data_214),
	.mem_107_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][107]~q ),
	.mem_107_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][107]~q ),
	.src_data_215(src_data_215),
	.mem_108_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][108]~q ),
	.mem_108_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][108]~q ),
	.src_data_216(src_data_216),
	.mem_109_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][109]~q ),
	.mem_109_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][109]~q ),
	.src_data_217(src_data_217),
	.mem_110_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][110]~q ),
	.mem_110_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][110]~q ),
	.src_data_218(src_data_218),
	.mem_111_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][111]~q ),
	.mem_111_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][111]~q ),
	.src_data_219(src_data_219),
	.mem_112_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][112]~q ),
	.mem_112_01(\onchip_sram_s2_agent_rsp_fifo|mem[0][112]~q ),
	.src_data_220(src_data_220));

Computer_System_Computer_System_mm_interconnect_0_rsp_demux_1 rsp_demux_001(
	.mem_66_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][66]~q ),
	.mem_68_0(\onchip_sram_s2_agent_rsp_fifo|mem[0][68]~q ),
	.src0_valid(\rsp_demux_001|src0_valid~0_combout ));

Computer_System_Computer_System_mm_interconnect_0_rsp_demux rsp_demux(
	.mem_68_0(\fifo_hps_to_fpga_in_agent_rsp_fifo|mem[0][68]~q ),
	.comb(\fifo_hps_to_fpga_in_agent|comb~0_combout ),
	.ShiftRight0(\fifo_hps_to_fpga_in_rsp_width_adapter|ShiftRight0~0_combout ),
	.always10(\fifo_hps_to_fpga_in_rsp_width_adapter|always10~0_combout ),
	.always101(\fifo_hps_to_fpga_in_rsp_width_adapter|always10~1_combout ),
	.src0_valid(\rsp_demux|src0_valid~0_combout ),
	.src1_valid(\rsp_demux|src1_valid~0_combout ));

endmodule

module Computer_System_altera_avalon_sc_fifo (
	clk,
	in_ready_hold,
	mem_31_0,
	reset)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	in_ready_hold;
output 	mem_31_0;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \mem[0][31] (
	.clk(clk),
	.d(in_ready_hold),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_31_0),
	.prn(vcc));
defparam \mem[0][31] .is_wysiwyg = "true";
defparam \mem[0][31] .power_up = "low";

endmodule

module Computer_System_altera_avalon_sc_fifo_1 (
	clk,
	out_valid_reg,
	mem_used_1,
	mem_68_0,
	mem_125_0,
	mem_used_0,
	comb,
	mem_122_0,
	mem_123_0,
	mem_124_0,
	mem_90_0,
	mem_91_0,
	ShiftRight0,
	mem_38_0,
	always10,
	mem_126_0,
	mem_39_0,
	always101,
	mem_101_0,
	mem_102_0,
	mem_103_0,
	mem_104_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	in_data_reg_68,
	nxt_uncomp_subburst_byte_cnt,
	reset,
	in_eop_reg,
	cp_ready,
	p1_ready,
	read,
	always102,
	in_data_reg_122,
	in_data_reg_123,
	in_data_reg_124,
	in_data_reg_90,
	in_data_reg_91,
	int_nxt_addr_reg_dly_2,
	mem_83_0,
	int_nxt_addr_reg_dly_3,
	mem_84_0,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	in_data_reg_104,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	out_burstwrap_reg_2,
	out_burstwrap_reg_3,
	mem_37_0,
	out_addr_reg_1,
	mem_82_0,
	mem_36_0,
	out_burstwrap_reg_1,
	out_addr_reg_0,
	mem_81_0,
	out_burstwrap_reg_0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	out_valid_reg;
output 	mem_used_1;
output 	mem_68_0;
output 	mem_125_0;
output 	mem_used_0;
input 	comb;
output 	mem_122_0;
output 	mem_123_0;
output 	mem_124_0;
output 	mem_90_0;
output 	mem_91_0;
input 	ShiftRight0;
output 	mem_38_0;
input 	always10;
output 	mem_126_0;
output 	mem_39_0;
input 	always101;
output 	mem_101_0;
output 	mem_102_0;
output 	mem_103_0;
output 	mem_104_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
input 	in_data_reg_68;
input 	nxt_uncomp_subburst_byte_cnt;
input 	reset;
input 	in_eop_reg;
input 	cp_ready;
input 	p1_ready;
output 	read;
input 	always102;
input 	in_data_reg_122;
input 	in_data_reg_123;
input 	in_data_reg_124;
input 	in_data_reg_90;
input 	in_data_reg_91;
input 	int_nxt_addr_reg_dly_2;
output 	mem_83_0;
input 	int_nxt_addr_reg_dly_3;
output 	mem_84_0;
input 	in_data_reg_101;
input 	in_data_reg_102;
input 	in_data_reg_103;
input 	in_data_reg_104;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
input 	out_burstwrap_reg_2;
input 	out_burstwrap_reg_3;
output 	mem_37_0;
input 	out_addr_reg_1;
output 	mem_82_0;
output 	mem_36_0;
input 	out_burstwrap_reg_1;
input 	out_addr_reg_0;
output 	mem_81_0;
input 	out_burstwrap_reg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][68]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][125]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][122]~q ;
wire \mem~2_combout ;
wire \mem[1][123]~q ;
wire \mem~3_combout ;
wire \mem[1][124]~q ;
wire \mem~4_combout ;
wire \mem[1][90]~q ;
wire \mem~5_combout ;
wire \mem[1][91]~q ;
wire \mem~6_combout ;
wire \mem[1][38]~q ;
wire \mem~7_combout ;
wire \mem[1][126]~q ;
wire \mem~8_combout ;
wire \mem[1][39]~q ;
wire \mem~9_combout ;
wire \mem[1][101]~q ;
wire \mem~10_combout ;
wire \mem[1][102]~q ;
wire \mem~11_combout ;
wire \mem[1][103]~q ;
wire \mem~12_combout ;
wire \mem[1][104]~q ;
wire \mem~13_combout ;
wire \mem[1][105]~q ;
wire \mem~14_combout ;
wire \mem[1][106]~q ;
wire \mem~15_combout ;
wire \mem[1][107]~q ;
wire \mem~16_combout ;
wire \mem[1][108]~q ;
wire \mem~17_combout ;
wire \mem[1][109]~q ;
wire \mem~18_combout ;
wire \mem[1][110]~q ;
wire \mem~19_combout ;
wire \mem[1][111]~q ;
wire \mem~20_combout ;
wire \mem[1][112]~q ;
wire \mem~21_combout ;
wire \mem[1][83]~q ;
wire \mem~22_combout ;
wire \mem[1][84]~q ;
wire \mem~23_combout ;
wire \mem[1][37]~q ;
wire \mem~24_combout ;
wire \mem[1][82]~q ;
wire \mem~25_combout ;
wire \mem[1][36]~q ;
wire \mem~26_combout ;
wire \mem[1][81]~q ;
wire \mem~27_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][125] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_125_0),
	.prn(vcc));
defparam \mem[0][125] .is_wysiwyg = "true";
defparam \mem[0][125] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][122] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_122_0),
	.prn(vcc));
defparam \mem[0][122] .is_wysiwyg = "true";
defparam \mem[0][122] .power_up = "low";

dffeas \mem[0][123] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_123_0),
	.prn(vcc));
defparam \mem[0][123] .is_wysiwyg = "true";
defparam \mem[0][123] .power_up = "low";

dffeas \mem[0][124] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_124_0),
	.prn(vcc));
defparam \mem[0][124] .is_wysiwyg = "true";
defparam \mem[0][124] .power_up = "low";

dffeas \mem[0][90] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_90_0),
	.prn(vcc));
defparam \mem[0][90] .is_wysiwyg = "true";
defparam \mem[0][90] .power_up = "low";

dffeas \mem[0][91] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_91_0),
	.prn(vcc));
defparam \mem[0][91] .is_wysiwyg = "true";
defparam \mem[0][91] .power_up = "low";

dffeas \mem[0][38] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_38_0),
	.prn(vcc));
defparam \mem[0][38] .is_wysiwyg = "true";
defparam \mem[0][38] .power_up = "low";

dffeas \mem[0][126] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_126_0),
	.prn(vcc));
defparam \mem[0][126] .is_wysiwyg = "true";
defparam \mem[0][126] .power_up = "low";

dffeas \mem[0][39] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_39_0),
	.prn(vcc));
defparam \mem[0][39] .is_wysiwyg = "true";
defparam \mem[0][39] .power_up = "low";

dffeas \mem[0][101] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_101_0),
	.prn(vcc));
defparam \mem[0][101] .is_wysiwyg = "true";
defparam \mem[0][101] .power_up = "low";

dffeas \mem[0][102] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_102_0),
	.prn(vcc));
defparam \mem[0][102] .is_wysiwyg = "true";
defparam \mem[0][102] .power_up = "low";

dffeas \mem[0][103] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_103_0),
	.prn(vcc));
defparam \mem[0][103] .is_wysiwyg = "true";
defparam \mem[0][103] .power_up = "low";

dffeas \mem[0][104] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_104_0),
	.prn(vcc));
defparam \mem[0][104] .is_wysiwyg = "true";
defparam \mem[0][104] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!ShiftRight0),
	.datac(!always10),
	.datad(!always101),
	.datae(!p1_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0051555500515555;
defparam \read~0 .shared_arith = "off";

dffeas \mem[0][83] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_83_0),
	.prn(vcc));
defparam \mem[0][83] .is_wysiwyg = "true";
defparam \mem[0][83] .power_up = "low";

dffeas \mem[0][84] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_84_0),
	.prn(vcc));
defparam \mem[0][84] .is_wysiwyg = "true";
defparam \mem[0][84] .power_up = "low";

dffeas \mem[0][37] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_37_0),
	.prn(vcc));
defparam \mem[0][37] .is_wysiwyg = "true";
defparam \mem[0][37] .power_up = "low";

dffeas \mem[0][82] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_82_0),
	.prn(vcc));
defparam \mem[0][82] .is_wysiwyg = "true";
defparam \mem[0][82] .power_up = "low";

dffeas \mem[0][36] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_36_0),
	.prn(vcc));
defparam \mem[0][36] .is_wysiwyg = "true";
defparam \mem[0][36] .power_up = "low";

dffeas \mem[0][81] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_81_0),
	.prn(vcc));
defparam \mem[0][81] .is_wysiwyg = "true";
defparam \mem[0][81] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!cp_ready),
	.datab(!in_data_reg_68),
	.datac(!nxt_uncomp_subburst_byte_cnt),
	.datad(!in_eop_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0001000100010001;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!read),
	.datad(!\write~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5035503550355035;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_68),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!read),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][125] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][125]~q ),
	.prn(vcc));
defparam \mem[1][125] .is_wysiwyg = "true";
defparam \mem[1][125] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!out_valid_reg),
	.datab(!mem_used_1),
	.datac(!in_data_reg_68),
	.datad(!in_eop_reg),
	.datae(!\mem[1][125]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h0004333700043337;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_125_0),
	.datac(!mem_used_0),
	.datad(!always102),
	.datae(!p1_ready),
	.dataf(!\write~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h0D0F0D0DFFFFFFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][122] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][122]~q ),
	.prn(vcc));
defparam \mem[1][122] .is_wysiwyg = "true";
defparam \mem[1][122] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][122]~q ),
	.datac(!in_data_reg_122),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][123] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][123]~q ),
	.prn(vcc));
defparam \mem[1][123] .is_wysiwyg = "true";
defparam \mem[1][123] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][123]~q ),
	.datac(!in_data_reg_123),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][124] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][124]~q ),
	.prn(vcc));
defparam \mem[1][124] .is_wysiwyg = "true";
defparam \mem[1][124] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][124]~q ),
	.datac(!in_data_reg_124),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][90] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][90]~q ),
	.prn(vcc));
defparam \mem[1][90] .is_wysiwyg = "true";
defparam \mem[1][90] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][90]~q ),
	.datac(!in_data_reg_90),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][91] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][91]~q ),
	.prn(vcc));
defparam \mem[1][91] .is_wysiwyg = "true";
defparam \mem[1][91] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][91]~q ),
	.datac(!in_data_reg_91),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][38] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][38]~q ),
	.prn(vcc));
defparam \mem[1][38] .is_wysiwyg = "true";
defparam \mem[1][38] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][38]~q ),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][126] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][126]~q ),
	.prn(vcc));
defparam \mem[1][126] .is_wysiwyg = "true";
defparam \mem[1][126] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!in_eop_reg),
	.datac(!\mem[1][126]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h2727272727272727;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][39] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][39]~q ),
	.prn(vcc));
defparam \mem[1][39] .is_wysiwyg = "true";
defparam \mem[1][39] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][39]~q ),
	.datac(!int_nxt_addr_reg_dly_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][101] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][101]~q ),
	.prn(vcc));
defparam \mem[1][101] .is_wysiwyg = "true";
defparam \mem[1][101] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][101]~q ),
	.datac(!in_data_reg_101),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][102] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][102]~q ),
	.prn(vcc));
defparam \mem[1][102] .is_wysiwyg = "true";
defparam \mem[1][102] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][102]~q ),
	.datac(!in_data_reg_102),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][103] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][103]~q ),
	.prn(vcc));
defparam \mem[1][103] .is_wysiwyg = "true";
defparam \mem[1][103] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][103]~q ),
	.datac(!in_data_reg_103),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][104] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][104]~q ),
	.prn(vcc));
defparam \mem[1][104] .is_wysiwyg = "true";
defparam \mem[1][104] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][104]~q ),
	.datac(!in_data_reg_104),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~20 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~21 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "off";
defparam \mem~21 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~21 .shared_arith = "off";

dffeas \mem[1][83] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][83]~q ),
	.prn(vcc));
defparam \mem[1][83] .is_wysiwyg = "true";
defparam \mem[1][83] .power_up = "low";

cyclonev_lcell_comb \mem~22 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][83]~q ),
	.datac(!out_burstwrap_reg_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~22 .extended_lut = "off";
defparam \mem~22 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~22 .shared_arith = "off";

dffeas \mem[1][84] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][84]~q ),
	.prn(vcc));
defparam \mem[1][84] .is_wysiwyg = "true";
defparam \mem[1][84] .power_up = "low";

cyclonev_lcell_comb \mem~23 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][84]~q ),
	.datac(!out_burstwrap_reg_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~23 .extended_lut = "off";
defparam \mem~23 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~23 .shared_arith = "off";

dffeas \mem[1][37] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][37]~q ),
	.prn(vcc));
defparam \mem[1][37] .is_wysiwyg = "true";
defparam \mem[1][37] .power_up = "low";

cyclonev_lcell_comb \mem~24 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][37]~q ),
	.datac(!out_addr_reg_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~24 .extended_lut = "off";
defparam \mem~24 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~24 .shared_arith = "off";

dffeas \mem[1][82] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][82]~q ),
	.prn(vcc));
defparam \mem[1][82] .is_wysiwyg = "true";
defparam \mem[1][82] .power_up = "low";

cyclonev_lcell_comb \mem~25 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][82]~q ),
	.datac(!out_burstwrap_reg_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~25 .extended_lut = "off";
defparam \mem~25 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~25 .shared_arith = "off";

dffeas \mem[1][36] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][36]~q ),
	.prn(vcc));
defparam \mem[1][36] .is_wysiwyg = "true";
defparam \mem[1][36] .power_up = "low";

cyclonev_lcell_comb \mem~26 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][36]~q ),
	.datac(!out_addr_reg_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~26 .extended_lut = "off";
defparam \mem~26 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~26 .shared_arith = "off";

dffeas \mem[1][81] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][81]~q ),
	.prn(vcc));
defparam \mem[1][81] .is_wysiwyg = "true";
defparam \mem[1][81] .power_up = "low";

cyclonev_lcell_comb \mem~27 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][81]~q ),
	.datac(!out_burstwrap_reg_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~27 .extended_lut = "off";
defparam \mem~27 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~27 .shared_arith = "off";

endmodule

module Computer_System_altera_avalon_sc_fifo_2 (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	clk,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_125_0,
	mem_used_01,
	out_valid,
	src_payload,
	always10,
	always4,
	mem_0_0,
	mem_1_0,
	mem_2_0,
	mem_3_0,
	mem_4_0,
	mem_5_0,
	mem_6_0,
	mem_7_0,
	mem_8_0,
	mem_9_0,
	mem_10_0,
	mem_11_0,
	mem_12_0,
	mem_13_0,
	mem_14_0,
	mem_15_0,
	mem_16_0,
	mem_17_0,
	mem_18_0,
	mem_19_0,
	mem_20_0,
	mem_21_0,
	mem_22_0,
	mem_23_0,
	mem_24_0,
	mem_25_0,
	mem_26_0,
	mem_27_0,
	mem_28_0,
	mem_29_0,
	mem_30_0,
	mem_31_0,
	out_data_1,
	out_data_4,
	out_data_6,
	out_data_8,
	out_data_13,
	out_data_17,
	out_data_20,
	out_data_22,
	out_data_24,
	out_data_29,
	reset,
	p1_ready)/* synthesis synthesis_greybox=0 */;
input 	q_b_0;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	q_b_8;
input 	q_b_9;
input 	q_b_10;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_20;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_24;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_28;
input 	q_b_29;
input 	q_b_30;
input 	q_b_31;
input 	clk;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_125_0;
input 	mem_used_01;
input 	out_valid;
input 	src_payload;
input 	always10;
output 	always4;
output 	mem_0_0;
output 	mem_1_0;
output 	mem_2_0;
output 	mem_3_0;
output 	mem_4_0;
output 	mem_5_0;
output 	mem_6_0;
output 	mem_7_0;
output 	mem_8_0;
output 	mem_9_0;
output 	mem_10_0;
output 	mem_11_0;
output 	mem_12_0;
output 	mem_13_0;
output 	mem_14_0;
output 	mem_15_0;
output 	mem_16_0;
output 	mem_17_0;
output 	mem_18_0;
output 	mem_19_0;
output 	mem_20_0;
output 	mem_21_0;
output 	mem_22_0;
output 	mem_23_0;
output 	mem_24_0;
output 	mem_25_0;
output 	mem_26_0;
output 	mem_27_0;
output 	mem_28_0;
output 	mem_29_0;
output 	mem_30_0;
output 	mem_31_0;
output 	out_data_1;
output 	out_data_4;
output 	out_data_6;
output 	out_data_8;
output 	out_data_13;
output 	out_data_17;
output 	out_data_20;
output 	out_data_22;
output 	out_data_24;
output 	out_data_29;
input 	reset;
input 	p1_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \read~1_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[1][8]~q ;
wire \mem~8_combout ;
wire \mem[1][9]~q ;
wire \mem~9_combout ;
wire \mem[1][10]~q ;
wire \mem~10_combout ;
wire \mem[1][11]~q ;
wire \mem~11_combout ;
wire \mem[1][12]~q ;
wire \mem~12_combout ;
wire \mem[1][13]~q ;
wire \mem~13_combout ;
wire \mem[1][14]~q ;
wire \mem~14_combout ;
wire \mem[1][15]~q ;
wire \mem~15_combout ;
wire \mem[1][16]~q ;
wire \mem~16_combout ;
wire \mem[1][17]~q ;
wire \mem~17_combout ;
wire \mem[1][18]~q ;
wire \mem~18_combout ;
wire \mem[1][19]~q ;
wire \mem~19_combout ;
wire \mem[1][20]~q ;
wire \mem~20_combout ;
wire \mem[1][21]~q ;
wire \mem~21_combout ;
wire \mem[1][22]~q ;
wire \mem~22_combout ;
wire \mem[1][23]~q ;
wire \mem~23_combout ;
wire \mem[1][24]~q ;
wire \mem~24_combout ;
wire \mem[1][25]~q ;
wire \mem~25_combout ;
wire \mem[1][26]~q ;
wire \mem~26_combout ;
wire \mem[1][27]~q ;
wire \mem~27_combout ;
wire \mem[1][28]~q ;
wire \mem~28_combout ;
wire \mem[1][29]~q ;
wire \mem~29_combout ;
wire \mem[1][30]~q ;
wire \mem~30_combout ;
wire \mem[1][31]~q ;
wire \mem~31_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \always4~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always4),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'h4444444444444444;
defparam \always4~0 .shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_8_0),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_9_0),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

dffeas \mem[0][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_10_0),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

dffeas \mem[0][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_11_0),
	.prn(vcc));
defparam \mem[0][11] .is_wysiwyg = "true";
defparam \mem[0][11] .power_up = "low";

dffeas \mem[0][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_12_0),
	.prn(vcc));
defparam \mem[0][12] .is_wysiwyg = "true";
defparam \mem[0][12] .power_up = "low";

dffeas \mem[0][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_13_0),
	.prn(vcc));
defparam \mem[0][13] .is_wysiwyg = "true";
defparam \mem[0][13] .power_up = "low";

dffeas \mem[0][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_14_0),
	.prn(vcc));
defparam \mem[0][14] .is_wysiwyg = "true";
defparam \mem[0][14] .power_up = "low";

dffeas \mem[0][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_15_0),
	.prn(vcc));
defparam \mem[0][15] .is_wysiwyg = "true";
defparam \mem[0][15] .power_up = "low";

dffeas \mem[0][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_16_0),
	.prn(vcc));
defparam \mem[0][16] .is_wysiwyg = "true";
defparam \mem[0][16] .power_up = "low";

dffeas \mem[0][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_17_0),
	.prn(vcc));
defparam \mem[0][17] .is_wysiwyg = "true";
defparam \mem[0][17] .power_up = "low";

dffeas \mem[0][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_18_0),
	.prn(vcc));
defparam \mem[0][18] .is_wysiwyg = "true";
defparam \mem[0][18] .power_up = "low";

dffeas \mem[0][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_19_0),
	.prn(vcc));
defparam \mem[0][19] .is_wysiwyg = "true";
defparam \mem[0][19] .power_up = "low";

dffeas \mem[0][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_20_0),
	.prn(vcc));
defparam \mem[0][20] .is_wysiwyg = "true";
defparam \mem[0][20] .power_up = "low";

dffeas \mem[0][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_21_0),
	.prn(vcc));
defparam \mem[0][21] .is_wysiwyg = "true";
defparam \mem[0][21] .power_up = "low";

dffeas \mem[0][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_22_0),
	.prn(vcc));
defparam \mem[0][22] .is_wysiwyg = "true";
defparam \mem[0][22] .power_up = "low";

dffeas \mem[0][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_23_0),
	.prn(vcc));
defparam \mem[0][23] .is_wysiwyg = "true";
defparam \mem[0][23] .power_up = "low";

dffeas \mem[0][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_24_0),
	.prn(vcc));
defparam \mem[0][24] .is_wysiwyg = "true";
defparam \mem[0][24] .power_up = "low";

dffeas \mem[0][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_25_0),
	.prn(vcc));
defparam \mem[0][25] .is_wysiwyg = "true";
defparam \mem[0][25] .power_up = "low";

dffeas \mem[0][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_26_0),
	.prn(vcc));
defparam \mem[0][26] .is_wysiwyg = "true";
defparam \mem[0][26] .power_up = "low";

dffeas \mem[0][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_27_0),
	.prn(vcc));
defparam \mem[0][27] .is_wysiwyg = "true";
defparam \mem[0][27] .power_up = "low";

dffeas \mem[0][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_28_0),
	.prn(vcc));
defparam \mem[0][28] .is_wysiwyg = "true";
defparam \mem[0][28] .power_up = "low";

dffeas \mem[0][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_29_0),
	.prn(vcc));
defparam \mem[0][29] .is_wysiwyg = "true";
defparam \mem[0][29] .power_up = "low";

dffeas \mem[0][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_30_0),
	.prn(vcc));
defparam \mem[0][30] .is_wysiwyg = "true";
defparam \mem[0][30] .power_up = "low";

dffeas \mem[0][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_31_0),
	.prn(vcc));
defparam \mem[0][31] .is_wysiwyg = "true";
defparam \mem[0][31] .power_up = "low";

cyclonev_lcell_comb \out_data[1]~0 (
	.dataa(!q_b_1),
	.datab(!always4),
	.datac(!mem_1_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[1]~0 .extended_lut = "off";
defparam \out_data[1]~0 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \out_data[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[4]~1 (
	.dataa(!q_b_4),
	.datab(!always4),
	.datac(!mem_4_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[4]~1 .extended_lut = "off";
defparam \out_data[4]~1 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \out_data[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[6]~2 (
	.dataa(!q_b_6),
	.datab(!always4),
	.datac(!mem_6_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[6]~2 .extended_lut = "off";
defparam \out_data[6]~2 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \out_data[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \out_data[8]~3 (
	.dataa(!q_b_8),
	.datab(!always4),
	.datac(!mem_8_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[8]~3 .extended_lut = "off";
defparam \out_data[8]~3 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \out_data[8]~3 .shared_arith = "off";

cyclonev_lcell_comb \out_data[13]~4 (
	.dataa(!q_b_13),
	.datab(!always4),
	.datac(!mem_13_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[13]~4 .extended_lut = "off";
defparam \out_data[13]~4 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \out_data[13]~4 .shared_arith = "off";

cyclonev_lcell_comb \out_data[17]~5 (
	.dataa(!q_b_17),
	.datab(!always4),
	.datac(!mem_17_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[17]~5 .extended_lut = "off";
defparam \out_data[17]~5 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \out_data[17]~5 .shared_arith = "off";

cyclonev_lcell_comb \out_data[20]~6 (
	.dataa(!q_b_20),
	.datab(!always4),
	.datac(!mem_20_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[20]~6 .extended_lut = "off";
defparam \out_data[20]~6 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \out_data[20]~6 .shared_arith = "off";

cyclonev_lcell_comb \out_data[22]~7 (
	.dataa(!q_b_22),
	.datab(!always4),
	.datac(!mem_22_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[22]~7 .extended_lut = "off";
defparam \out_data[22]~7 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \out_data[22]~7 .shared_arith = "off";

cyclonev_lcell_comb \out_data[24]~8 (
	.dataa(!q_b_24),
	.datab(!always4),
	.datac(!mem_24_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[24]~8 .extended_lut = "off";
defparam \out_data[24]~8 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \out_data[24]~8 .shared_arith = "off";

cyclonev_lcell_comb \out_data[29]~9 (
	.dataa(!q_b_29),
	.datab(!always4),
	.datac(!mem_29_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[29]~9 .extended_lut = "off";
defparam \out_data[29]~9 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \out_data[29]~9 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_125_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h888F888F888F888F;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \read~1 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!p1_ready),
	.datae(!\read~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~1 .extended_lut = "off";
defparam \read~1 .lut_mask = 64'h5DFF00005DFF0000;
defparam \read~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!q_b_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!out_valid),
	.datac(!src_payload),
	.datad(!always10),
	.datae(!p1_ready),
	.dataf(!\read~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBFBFFFFAAAAAAAA;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!q_b_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!q_b_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!q_b_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!q_b_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!q_b_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!q_b_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!q_b_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!q_b_8),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!q_b_9),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h4747474747474747;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!q_b_10),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h4747474747474747;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][11]~q ),
	.prn(vcc));
defparam \mem[1][11] .is_wysiwyg = "true";
defparam \mem[1][11] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!q_b_11),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h4747474747474747;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][12]~q ),
	.prn(vcc));
defparam \mem[1][12] .is_wysiwyg = "true";
defparam \mem[1][12] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!q_b_12),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h4747474747474747;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][13]~q ),
	.prn(vcc));
defparam \mem[1][13] .is_wysiwyg = "true";
defparam \mem[1][13] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!q_b_13),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h4747474747474747;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][14]~q ),
	.prn(vcc));
defparam \mem[1][14] .is_wysiwyg = "true";
defparam \mem[1][14] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!q_b_14),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h4747474747474747;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][15]~q ),
	.prn(vcc));
defparam \mem[1][15] .is_wysiwyg = "true";
defparam \mem[1][15] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!q_b_15),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h4747474747474747;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][16]~q ),
	.prn(vcc));
defparam \mem[1][16] .is_wysiwyg = "true";
defparam \mem[1][16] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!q_b_16),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][16]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h4747474747474747;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][17]~q ),
	.prn(vcc));
defparam \mem[1][17] .is_wysiwyg = "true";
defparam \mem[1][17] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!q_b_17),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h4747474747474747;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][18]~q ),
	.prn(vcc));
defparam \mem[1][18] .is_wysiwyg = "true";
defparam \mem[1][18] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!q_b_18),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h4747474747474747;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][19]~q ),
	.prn(vcc));
defparam \mem[1][19] .is_wysiwyg = "true";
defparam \mem[1][19] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!q_b_19),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h4747474747474747;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[1][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][20]~q ),
	.prn(vcc));
defparam \mem[1][20] .is_wysiwyg = "true";
defparam \mem[1][20] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!q_b_20),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h4747474747474747;
defparam \mem~20 .shared_arith = "off";

dffeas \mem[1][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][21]~q ),
	.prn(vcc));
defparam \mem[1][21] .is_wysiwyg = "true";
defparam \mem[1][21] .power_up = "low";

cyclonev_lcell_comb \mem~21 (
	.dataa(!q_b_21),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "off";
defparam \mem~21 .lut_mask = 64'h4747474747474747;
defparam \mem~21 .shared_arith = "off";

dffeas \mem[1][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][22]~q ),
	.prn(vcc));
defparam \mem[1][22] .is_wysiwyg = "true";
defparam \mem[1][22] .power_up = "low";

cyclonev_lcell_comb \mem~22 (
	.dataa(!q_b_22),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~22 .extended_lut = "off";
defparam \mem~22 .lut_mask = 64'h4747474747474747;
defparam \mem~22 .shared_arith = "off";

dffeas \mem[1][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][23]~q ),
	.prn(vcc));
defparam \mem[1][23] .is_wysiwyg = "true";
defparam \mem[1][23] .power_up = "low";

cyclonev_lcell_comb \mem~23 (
	.dataa(!q_b_23),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~23 .extended_lut = "off";
defparam \mem~23 .lut_mask = 64'h4747474747474747;
defparam \mem~23 .shared_arith = "off";

dffeas \mem[1][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][24]~q ),
	.prn(vcc));
defparam \mem[1][24] .is_wysiwyg = "true";
defparam \mem[1][24] .power_up = "low";

cyclonev_lcell_comb \mem~24 (
	.dataa(!q_b_24),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~24 .extended_lut = "off";
defparam \mem~24 .lut_mask = 64'h4747474747474747;
defparam \mem~24 .shared_arith = "off";

dffeas \mem[1][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][25]~q ),
	.prn(vcc));
defparam \mem[1][25] .is_wysiwyg = "true";
defparam \mem[1][25] .power_up = "low";

cyclonev_lcell_comb \mem~25 (
	.dataa(!q_b_25),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~25 .extended_lut = "off";
defparam \mem~25 .lut_mask = 64'h4747474747474747;
defparam \mem~25 .shared_arith = "off";

dffeas \mem[1][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][26]~q ),
	.prn(vcc));
defparam \mem[1][26] .is_wysiwyg = "true";
defparam \mem[1][26] .power_up = "low";

cyclonev_lcell_comb \mem~26 (
	.dataa(!q_b_26),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~26 .extended_lut = "off";
defparam \mem~26 .lut_mask = 64'h4747474747474747;
defparam \mem~26 .shared_arith = "off";

dffeas \mem[1][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][27]~q ),
	.prn(vcc));
defparam \mem[1][27] .is_wysiwyg = "true";
defparam \mem[1][27] .power_up = "low";

cyclonev_lcell_comb \mem~27 (
	.dataa(!q_b_27),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~27 .extended_lut = "off";
defparam \mem~27 .lut_mask = 64'h4747474747474747;
defparam \mem~27 .shared_arith = "off";

dffeas \mem[1][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][28]~q ),
	.prn(vcc));
defparam \mem[1][28] .is_wysiwyg = "true";
defparam \mem[1][28] .power_up = "low";

cyclonev_lcell_comb \mem~28 (
	.dataa(!q_b_28),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~28 .extended_lut = "off";
defparam \mem~28 .lut_mask = 64'h4747474747474747;
defparam \mem~28 .shared_arith = "off";

dffeas \mem[1][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][29]~q ),
	.prn(vcc));
defparam \mem[1][29] .is_wysiwyg = "true";
defparam \mem[1][29] .power_up = "low";

cyclonev_lcell_comb \mem~29 (
	.dataa(!q_b_29),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~29 .extended_lut = "off";
defparam \mem~29 .lut_mask = 64'h4747474747474747;
defparam \mem~29 .shared_arith = "off";

dffeas \mem[1][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][30]~q ),
	.prn(vcc));
defparam \mem[1][30] .is_wysiwyg = "true";
defparam \mem[1][30] .power_up = "low";

cyclonev_lcell_comb \mem~30 (
	.dataa(!q_b_30),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~30 .extended_lut = "off";
defparam \mem~30 .lut_mask = 64'h4747474747474747;
defparam \mem~30 .shared_arith = "off";

dffeas \mem[1][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][31]~q ),
	.prn(vcc));
defparam \mem[1][31] .is_wysiwyg = "true";
defparam \mem[1][31] .power_up = "low";

cyclonev_lcell_comb \mem~31 (
	.dataa(!q_b_31),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~31 .extended_lut = "off";
defparam \mem~31 .lut_mask = 64'h4747474747474747;
defparam \mem~31 .shared_arith = "off";

endmodule

module Computer_System_altera_avalon_sc_fifo_3 (
	clk,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_7,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_8,
	out_uncomp_byte_cnt_reg_5,
	out_burstwrap_reg_2,
	out_burstwrap_reg_3,
	out_addr_reg_1,
	out_burstwrap_reg_1,
	out_addr_reg_0,
	out_burstwrap_reg_0,
	stateST_COMP_TRANS,
	in_data_reg_91,
	in_data_reg_90,
	mem_used_1,
	cp_ready,
	in_eop_reg,
	new_burst_reg,
	in_bytecount_reg_zero,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	mem_125_0,
	mem_used_0,
	out_valid,
	comb,
	mem_126_0,
	mem_66_0,
	mem_80_0,
	mem_79_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	mem_38_0,
	mem_122_0,
	mem_123_0,
	mem_91_0,
	mem_124_0,
	mem_90_0,
	mem_39_0,
	always10,
	mem_68_0,
	mem_101_0,
	mem_102_0,
	mem_103_0,
	mem_104_0,
	mem_105_0,
	mem_106_0,
	mem_107_0,
	mem_108_0,
	mem_109_0,
	mem_110_0,
	mem_111_0,
	mem_112_0,
	in_data_reg_68,
	reset,
	nxt_out_eop,
	in_data_reg_69,
	last_packet_beat,
	p1_ready,
	cp_ready1,
	out_byte_cnt_reg_2,
	WideOr0,
	always101,
	mem_83_0,
	in_data_reg_122,
	in_data_reg_123,
	in_data_reg_124,
	mem_84_0,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	in_data_reg_104,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	mem_37_0,
	mem_82_0,
	mem_36_0,
	mem_81_0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	int_nxt_addr_reg_dly_2;
input 	int_nxt_addr_reg_dly_3;
input 	out_uncomp_byte_cnt_reg_6;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_7;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_8;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_burstwrap_reg_2;
input 	out_burstwrap_reg_3;
input 	out_addr_reg_1;
input 	out_burstwrap_reg_1;
input 	out_addr_reg_0;
input 	out_burstwrap_reg_0;
input 	stateST_COMP_TRANS;
input 	in_data_reg_91;
input 	in_data_reg_90;
output 	mem_used_1;
input 	cp_ready;
input 	in_eop_reg;
input 	new_burst_reg;
input 	in_bytecount_reg_zero;
input 	out_valid_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_125_0;
output 	mem_used_0;
input 	out_valid;
input 	comb;
output 	mem_126_0;
output 	mem_66_0;
output 	mem_80_0;
output 	mem_79_0;
output 	mem_78_0;
output 	mem_77_0;
output 	mem_76_0;
output 	mem_75_0;
output 	mem_74_0;
output 	mem_38_0;
output 	mem_122_0;
output 	mem_123_0;
output 	mem_91_0;
output 	mem_124_0;
output 	mem_90_0;
output 	mem_39_0;
input 	always10;
output 	mem_68_0;
output 	mem_101_0;
output 	mem_102_0;
output 	mem_103_0;
output 	mem_104_0;
output 	mem_105_0;
output 	mem_106_0;
output 	mem_107_0;
output 	mem_108_0;
output 	mem_109_0;
output 	mem_110_0;
output 	mem_111_0;
output 	mem_112_0;
input 	in_data_reg_68;
input 	reset;
input 	nxt_out_eop;
input 	in_data_reg_69;
input 	last_packet_beat;
input 	p1_ready;
input 	cp_ready1;
input 	out_byte_cnt_reg_2;
input 	WideOr0;
input 	always101;
output 	mem_83_0;
input 	in_data_reg_122;
input 	in_data_reg_123;
input 	in_data_reg_124;
output 	mem_84_0;
input 	in_data_reg_101;
input 	in_data_reg_102;
input 	in_data_reg_103;
input 	in_data_reg_104;
input 	in_data_reg_105;
input 	in_data_reg_106;
input 	in_data_reg_107;
input 	in_data_reg_108;
input 	in_data_reg_109;
input 	in_data_reg_110;
input 	in_data_reg_111;
input 	in_data_reg_112;
output 	mem_37_0;
output 	mem_82_0;
output 	mem_36_0;
output 	mem_81_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \read~0_combout ;
wire \write~1_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][125]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][126]~q ;
wire \mem~1_combout ;
wire \mem[1][69]~q ;
wire \mem~2_combout ;
wire \mem[1][80]~q ;
wire \mem~3_combout ;
wire \mem[1][79]~q ;
wire \mem~4_combout ;
wire \mem[1][78]~q ;
wire \mem~5_combout ;
wire \mem[1][77]~q ;
wire \mem~6_combout ;
wire \mem[1][76]~q ;
wire \mem~7_combout ;
wire \mem[1][75]~q ;
wire \mem~8_combout ;
wire \mem[1][74]~q ;
wire \mem~9_combout ;
wire \mem[1][38]~q ;
wire \mem~10_combout ;
wire \mem[1][122]~q ;
wire \mem~11_combout ;
wire \mem[1][123]~q ;
wire \mem~12_combout ;
wire \mem[1][91]~q ;
wire \mem~13_combout ;
wire \mem[1][124]~q ;
wire \mem~14_combout ;
wire \mem[1][90]~q ;
wire \mem~15_combout ;
wire \mem[1][39]~q ;
wire \mem~16_combout ;
wire \mem[1][68]~q ;
wire \mem~17_combout ;
wire \mem[1][101]~q ;
wire \mem~18_combout ;
wire \mem[1][102]~q ;
wire \mem~19_combout ;
wire \mem[1][103]~q ;
wire \mem~20_combout ;
wire \mem[1][104]~q ;
wire \mem~21_combout ;
wire \mem[1][105]~q ;
wire \mem~22_combout ;
wire \mem[1][106]~q ;
wire \mem~23_combout ;
wire \mem[1][107]~q ;
wire \mem~24_combout ;
wire \mem[1][108]~q ;
wire \mem~25_combout ;
wire \mem[1][109]~q ;
wire \mem~26_combout ;
wire \mem[1][110]~q ;
wire \mem~27_combout ;
wire \mem[1][111]~q ;
wire \mem~28_combout ;
wire \mem[1][112]~q ;
wire \mem~29_combout ;
wire \mem[1][83]~q ;
wire \mem~30_combout ;
wire \mem[1][84]~q ;
wire \mem~31_combout ;
wire \mem[1][37]~q ;
wire \mem~32_combout ;
wire \mem[1][82]~q ;
wire \mem~33_combout ;
wire \mem[1][36]~q ;
wire \mem~34_combout ;
wire \mem[1][81]~q ;
wire \mem~35_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][125] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_125_0),
	.prn(vcc));
defparam \mem[0][125] .is_wysiwyg = "true";
defparam \mem[0][125] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][126] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_126_0),
	.prn(vcc));
defparam \mem[0][126] .is_wysiwyg = "true";
defparam \mem[0][126] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][80] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_80_0),
	.prn(vcc));
defparam \mem[0][80] .is_wysiwyg = "true";
defparam \mem[0][80] .power_up = "low";

dffeas \mem[0][79] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_79_0),
	.prn(vcc));
defparam \mem[0][79] .is_wysiwyg = "true";
defparam \mem[0][79] .power_up = "low";

dffeas \mem[0][78] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_78_0),
	.prn(vcc));
defparam \mem[0][78] .is_wysiwyg = "true";
defparam \mem[0][78] .power_up = "low";

dffeas \mem[0][77] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_77_0),
	.prn(vcc));
defparam \mem[0][77] .is_wysiwyg = "true";
defparam \mem[0][77] .power_up = "low";

dffeas \mem[0][76] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_76_0),
	.prn(vcc));
defparam \mem[0][76] .is_wysiwyg = "true";
defparam \mem[0][76] .power_up = "low";

dffeas \mem[0][75] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_75_0),
	.prn(vcc));
defparam \mem[0][75] .is_wysiwyg = "true";
defparam \mem[0][75] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][38] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_38_0),
	.prn(vcc));
defparam \mem[0][38] .is_wysiwyg = "true";
defparam \mem[0][38] .power_up = "low";

dffeas \mem[0][122] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_122_0),
	.prn(vcc));
defparam \mem[0][122] .is_wysiwyg = "true";
defparam \mem[0][122] .power_up = "low";

dffeas \mem[0][123] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_123_0),
	.prn(vcc));
defparam \mem[0][123] .is_wysiwyg = "true";
defparam \mem[0][123] .power_up = "low";

dffeas \mem[0][91] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_91_0),
	.prn(vcc));
defparam \mem[0][91] .is_wysiwyg = "true";
defparam \mem[0][91] .power_up = "low";

dffeas \mem[0][124] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_124_0),
	.prn(vcc));
defparam \mem[0][124] .is_wysiwyg = "true";
defparam \mem[0][124] .power_up = "low";

dffeas \mem[0][90] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_90_0),
	.prn(vcc));
defparam \mem[0][90] .is_wysiwyg = "true";
defparam \mem[0][90] .power_up = "low";

dffeas \mem[0][39] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_39_0),
	.prn(vcc));
defparam \mem[0][39] .is_wysiwyg = "true";
defparam \mem[0][39] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][101] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_101_0),
	.prn(vcc));
defparam \mem[0][101] .is_wysiwyg = "true";
defparam \mem[0][101] .power_up = "low";

dffeas \mem[0][102] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_102_0),
	.prn(vcc));
defparam \mem[0][102] .is_wysiwyg = "true";
defparam \mem[0][102] .power_up = "low";

dffeas \mem[0][103] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_103_0),
	.prn(vcc));
defparam \mem[0][103] .is_wysiwyg = "true";
defparam \mem[0][103] .power_up = "low";

dffeas \mem[0][104] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_104_0),
	.prn(vcc));
defparam \mem[0][104] .is_wysiwyg = "true";
defparam \mem[0][104] .power_up = "low";

dffeas \mem[0][105] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_105_0),
	.prn(vcc));
defparam \mem[0][105] .is_wysiwyg = "true";
defparam \mem[0][105] .power_up = "low";

dffeas \mem[0][106] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_106_0),
	.prn(vcc));
defparam \mem[0][106] .is_wysiwyg = "true";
defparam \mem[0][106] .power_up = "low";

dffeas \mem[0][107] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_107_0),
	.prn(vcc));
defparam \mem[0][107] .is_wysiwyg = "true";
defparam \mem[0][107] .power_up = "low";

dffeas \mem[0][108] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_108_0),
	.prn(vcc));
defparam \mem[0][108] .is_wysiwyg = "true";
defparam \mem[0][108] .power_up = "low";

dffeas \mem[0][109] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_109_0),
	.prn(vcc));
defparam \mem[0][109] .is_wysiwyg = "true";
defparam \mem[0][109] .power_up = "low";

dffeas \mem[0][110] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_110_0),
	.prn(vcc));
defparam \mem[0][110] .is_wysiwyg = "true";
defparam \mem[0][110] .power_up = "low";

dffeas \mem[0][111] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_111_0),
	.prn(vcc));
defparam \mem[0][111] .is_wysiwyg = "true";
defparam \mem[0][111] .power_up = "low";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem[0][83] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_83_0),
	.prn(vcc));
defparam \mem[0][83] .is_wysiwyg = "true";
defparam \mem[0][83] .power_up = "low";

dffeas \mem[0][84] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_84_0),
	.prn(vcc));
defparam \mem[0][84] .is_wysiwyg = "true";
defparam \mem[0][84] .power_up = "low";

dffeas \mem[0][37] (
	.clk(clk),
	.d(\mem~32_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_37_0),
	.prn(vcc));
defparam \mem[0][37] .is_wysiwyg = "true";
defparam \mem[0][37] .power_up = "low";

dffeas \mem[0][82] (
	.clk(clk),
	.d(\mem~33_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_82_0),
	.prn(vcc));
defparam \mem[0][82] .is_wysiwyg = "true";
defparam \mem[0][82] .power_up = "low";

dffeas \mem[0][36] (
	.clk(clk),
	.d(\mem~34_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_36_0),
	.prn(vcc));
defparam \mem[0][36] .is_wysiwyg = "true";
defparam \mem[0][36] .power_up = "low";

dffeas \mem[0][81] (
	.clk(clk),
	.d(\mem~35_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_81_0),
	.prn(vcc));
defparam \mem[0][81] .is_wysiwyg = "true";
defparam \mem[0][81] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!cp_ready),
	.datac(!in_eop_reg),
	.datad(!new_burst_reg),
	.datae(!in_bytecount_reg_zero),
	.dataf(!in_data_reg_68),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h000000000A1B4E5F;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!out_valid),
	.datac(!mem_126_0),
	.datad(!last_packet_beat),
	.datae(!always10),
	.dataf(!p1_ready),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0011005100550055;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!out_valid_reg),
	.datab(!cp_ready1),
	.datac(!mem_used_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h1010101010101010;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!in_data_reg_69),
	.datad(!\write~0_combout ),
	.datae(!\read~0_combout ),
	.dataf(!\write~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5555000053330555;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][125] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][125]~q ),
	.prn(vcc));
defparam \mem[1][125] .is_wysiwyg = "true";
defparam \mem[1][125] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!out_valid_reg),
	.datab(!WideOr0),
	.datac(!mem_used_1),
	.datad(!in_data_reg_69),
	.datae(!\write~0_combout ),
	.dataf(!\mem[1][125]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h001050500F1F5F5F;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!comb),
	.datac(!out_valid),
	.datad(!last_packet_beat),
	.datae(!always101),
	.dataf(!p1_ready),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hAABBAAABAABBAABB;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!in_data_reg_69),
	.datad(!\write~0_combout ),
	.datae(!\read~0_combout ),
	.dataf(!\write~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h333311113FFF1FFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][126] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][126]~q ),
	.prn(vcc));
defparam \mem[1][126] .is_wysiwyg = "true";
defparam \mem[1][126] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][126]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_69),
	.datac(!\mem[1][69]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][80] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][80]~q ),
	.prn(vcc));
defparam \mem[1][80] .is_wysiwyg = "true";
defparam \mem[1][80] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_8),
	.datad(!\mem[1][80]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][79] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][79]~q ),
	.prn(vcc));
defparam \mem[1][79] .is_wysiwyg = "true";
defparam \mem[1][79] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_7),
	.datad(!\mem[1][79]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][78] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][78]~q ),
	.prn(vcc));
defparam \mem[1][78] .is_wysiwyg = "true";
defparam \mem[1][78] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][77] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][77]~q ),
	.prn(vcc));
defparam \mem[1][77] .is_wysiwyg = "true";
defparam \mem[1][77] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][76] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][76]~q ),
	.prn(vcc));
defparam \mem[1][76] .is_wysiwyg = "true";
defparam \mem[1][76] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h0257025702570257;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][75] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][75]~q ),
	.prn(vcc));
defparam \mem[1][75] .is_wysiwyg = "true";
defparam \mem[1][75] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h0257025702570257;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][74]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][38] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][38]~q ),
	.prn(vcc));
defparam \mem[1][38] .is_wysiwyg = "true";
defparam \mem[1][38] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!\mem[1][38]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h2727272727272727;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][122] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][122]~q ),
	.prn(vcc));
defparam \mem[1][122] .is_wysiwyg = "true";
defparam \mem[1][122] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][122]~q ),
	.datac(!in_data_reg_122),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][123] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][123]~q ),
	.prn(vcc));
defparam \mem[1][123] .is_wysiwyg = "true";
defparam \mem[1][123] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][123]~q ),
	.datac(!in_data_reg_123),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][91] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][91]~q ),
	.prn(vcc));
defparam \mem[1][91] .is_wysiwyg = "true";
defparam \mem[1][91] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!in_data_reg_91),
	.datab(!mem_used_1),
	.datac(!\mem[1][91]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h4747474747474747;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][124] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][124]~q ),
	.prn(vcc));
defparam \mem[1][124] .is_wysiwyg = "true";
defparam \mem[1][124] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][124]~q ),
	.datac(!in_data_reg_124),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][90] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][90]~q ),
	.prn(vcc));
defparam \mem[1][90] .is_wysiwyg = "true";
defparam \mem[1][90] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!in_data_reg_90),
	.datab(!mem_used_1),
	.datac(!\mem[1][90]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h4747474747474747;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][39] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][39]~q ),
	.prn(vcc));
defparam \mem[1][39] .is_wysiwyg = "true";
defparam \mem[1][39] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!\mem[1][39]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h2727272727272727;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_68),
	.datac(!\mem[1][68]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h2727272727272727;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][101] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][101]~q ),
	.prn(vcc));
defparam \mem[1][101] .is_wysiwyg = "true";
defparam \mem[1][101] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][101]~q ),
	.datac(!in_data_reg_101),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][102] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][102]~q ),
	.prn(vcc));
defparam \mem[1][102] .is_wysiwyg = "true";
defparam \mem[1][102] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][102]~q ),
	.datac(!in_data_reg_102),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[1][103] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][103]~q ),
	.prn(vcc));
defparam \mem[1][103] .is_wysiwyg = "true";
defparam \mem[1][103] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][103]~q ),
	.datac(!in_data_reg_103),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~20 .shared_arith = "off";

dffeas \mem[1][104] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][104]~q ),
	.prn(vcc));
defparam \mem[1][104] .is_wysiwyg = "true";
defparam \mem[1][104] .power_up = "low";

cyclonev_lcell_comb \mem~21 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][104]~q ),
	.datac(!in_data_reg_104),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "off";
defparam \mem~21 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~21 .shared_arith = "off";

dffeas \mem[1][105] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][105]~q ),
	.prn(vcc));
defparam \mem[1][105] .is_wysiwyg = "true";
defparam \mem[1][105] .power_up = "low";

cyclonev_lcell_comb \mem~22 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][105]~q ),
	.datac(!in_data_reg_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~22 .extended_lut = "off";
defparam \mem~22 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~22 .shared_arith = "off";

dffeas \mem[1][106] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][106]~q ),
	.prn(vcc));
defparam \mem[1][106] .is_wysiwyg = "true";
defparam \mem[1][106] .power_up = "low";

cyclonev_lcell_comb \mem~23 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][106]~q ),
	.datac(!in_data_reg_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~23 .extended_lut = "off";
defparam \mem~23 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~23 .shared_arith = "off";

dffeas \mem[1][107] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][107]~q ),
	.prn(vcc));
defparam \mem[1][107] .is_wysiwyg = "true";
defparam \mem[1][107] .power_up = "low";

cyclonev_lcell_comb \mem~24 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][107]~q ),
	.datac(!in_data_reg_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~24 .extended_lut = "off";
defparam \mem~24 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~24 .shared_arith = "off";

dffeas \mem[1][108] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][108]~q ),
	.prn(vcc));
defparam \mem[1][108] .is_wysiwyg = "true";
defparam \mem[1][108] .power_up = "low";

cyclonev_lcell_comb \mem~25 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][108]~q ),
	.datac(!in_data_reg_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~25 .extended_lut = "off";
defparam \mem~25 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~25 .shared_arith = "off";

dffeas \mem[1][109] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][109]~q ),
	.prn(vcc));
defparam \mem[1][109] .is_wysiwyg = "true";
defparam \mem[1][109] .power_up = "low";

cyclonev_lcell_comb \mem~26 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][109]~q ),
	.datac(!in_data_reg_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~26 .extended_lut = "off";
defparam \mem~26 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~26 .shared_arith = "off";

dffeas \mem[1][110] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][110]~q ),
	.prn(vcc));
defparam \mem[1][110] .is_wysiwyg = "true";
defparam \mem[1][110] .power_up = "low";

cyclonev_lcell_comb \mem~27 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][110]~q ),
	.datac(!in_data_reg_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~27 .extended_lut = "off";
defparam \mem~27 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~27 .shared_arith = "off";

dffeas \mem[1][111] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][111]~q ),
	.prn(vcc));
defparam \mem[1][111] .is_wysiwyg = "true";
defparam \mem[1][111] .power_up = "low";

cyclonev_lcell_comb \mem~28 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][111]~q ),
	.datac(!in_data_reg_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~28 .extended_lut = "off";
defparam \mem~28 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~28 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~29 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][112]~q ),
	.datac(!in_data_reg_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~29 .extended_lut = "off";
defparam \mem~29 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~29 .shared_arith = "off";

dffeas \mem[1][83] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][83]~q ),
	.prn(vcc));
defparam \mem[1][83] .is_wysiwyg = "true";
defparam \mem[1][83] .power_up = "low";

cyclonev_lcell_comb \mem~30 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][83]~q ),
	.datac(!out_burstwrap_reg_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~30 .extended_lut = "off";
defparam \mem~30 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~30 .shared_arith = "off";

dffeas \mem[1][84] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][84]~q ),
	.prn(vcc));
defparam \mem[1][84] .is_wysiwyg = "true";
defparam \mem[1][84] .power_up = "low";

cyclonev_lcell_comb \mem~31 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][84]~q ),
	.datac(!out_burstwrap_reg_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~31 .extended_lut = "off";
defparam \mem~31 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~31 .shared_arith = "off";

dffeas \mem[1][37] (
	.clk(clk),
	.d(\mem~32_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][37]~q ),
	.prn(vcc));
defparam \mem[1][37] .is_wysiwyg = "true";
defparam \mem[1][37] .power_up = "low";

cyclonev_lcell_comb \mem~32 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][37]~q ),
	.datac(!out_addr_reg_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~32 .extended_lut = "off";
defparam \mem~32 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~32 .shared_arith = "off";

dffeas \mem[1][82] (
	.clk(clk),
	.d(\mem~33_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][82]~q ),
	.prn(vcc));
defparam \mem[1][82] .is_wysiwyg = "true";
defparam \mem[1][82] .power_up = "low";

cyclonev_lcell_comb \mem~33 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][82]~q ),
	.datac(!out_burstwrap_reg_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~33 .extended_lut = "off";
defparam \mem~33 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~33 .shared_arith = "off";

dffeas \mem[1][36] (
	.clk(clk),
	.d(\mem~34_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][36]~q ),
	.prn(vcc));
defparam \mem[1][36] .is_wysiwyg = "true";
defparam \mem[1][36] .power_up = "low";

cyclonev_lcell_comb \mem~34 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][36]~q ),
	.datac(!out_addr_reg_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~34 .extended_lut = "off";
defparam \mem~34 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~34 .shared_arith = "off";

dffeas \mem[1][81] (
	.clk(clk),
	.d(\mem~35_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][81]~q ),
	.prn(vcc));
defparam \mem[1][81] .is_wysiwyg = "true";
defparam \mem[1][81] .power_up = "low";

cyclonev_lcell_comb \mem~35 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][81]~q ),
	.datac(!out_burstwrap_reg_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~35 .extended_lut = "off";
defparam \mem~35 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~35 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_axi_master_ni (
	h2f_WLAST_0,
	h2f_ARLEN_0,
	h2f_ARLEN_1,
	h2f_ARLEN_2,
	h2f_ARLEN_3,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWADDR_0,
	h2f_AWADDR_1,
	h2f_AWADDR_2,
	h2f_AWADDR_3,
	h2f_AWADDR_4,
	h2f_AWADDR_5,
	h2f_AWADDR_6,
	h2f_AWADDR_7,
	h2f_AWADDR_8,
	h2f_AWADDR_9,
	h2f_AWADDR_10,
	h2f_AWADDR_11,
	h2f_AWADDR_12,
	h2f_AWADDR_13,
	h2f_AWADDR_14,
	h2f_AWADDR_15,
	h2f_AWADDR_16,
	h2f_AWADDR_17,
	h2f_AWADDR_18,
	h2f_AWADDR_19,
	h2f_AWADDR_20,
	h2f_AWADDR_21,
	h2f_AWADDR_22,
	h2f_AWADDR_23,
	h2f_AWADDR_24,
	h2f_AWADDR_25,
	h2f_AWADDR_26,
	h2f_AWADDR_27,
	h2f_AWBURST_0,
	h2f_AWBURST_1,
	h2f_AWLEN_0,
	h2f_AWLEN_1,
	h2f_AWLEN_2,
	h2f_AWLEN_3,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	outclk_wire_0,
	address_burst_24,
	address_burst_25,
	address_burst_23,
	address_burst_13,
	address_burst_21,
	address_burst_22,
	address_burst_19,
	address_burst_20,
	address_burst_15,
	address_burst_16,
	address_burst_17,
	address_burst_18,
	address_burst_26,
	address_burst_27,
	address_burst_12,
	address_burst_14,
	address_burst_10,
	address_burst_11,
	address_burst_9,
	address_burst_8,
	Add4,
	Add5,
	Add41,
	Add51,
	Add42,
	Add52,
	Add43,
	Add53,
	Add44,
	Add54,
	Add55,
	Add45,
	Add56,
	Add46,
	Add47,
	Add57,
	Add48,
	Add58,
	in_ready,
	nxt_in_ready,
	sop_enable1,
	address_burst_7,
	address_burst_6,
	address_burst_2,
	address_burst_3,
	address_burst_4,
	address_burst_5,
	sink_ready,
	sink_ready1,
	cmd_sink_ready,
	last_cycle,
	awready,
	last_cycle1,
	wready,
	LessThan11,
	Add3,
	log2ceil,
	address_burst_1,
	LessThan10,
	Add31,
	address_burst_0,
	out_data_2,
	out_data_3,
	burst_bytecount_4,
	burst_bytecount_6,
	burst_bytecount_5,
	burst_bytecount_7,
	Add0,
	Add2,
	Add01,
	Add21,
	Add22,
	write_cp_data_188,
	write_cp_data_187,
	altera_reset_synchronizer_int_chain_out,
	out_data_7,
	Add1,
	out_data_9,
	out_data_6,
	LessThan16,
	out_data_8,
	LessThan12,
	Selector26,
	out_data_4,
	LessThan14,
	out_data_5,
	LessThan15,
	LessThan2,
	Add32,
	Selector7,
	out_data_1,
	Decoder0,
	Selector8,
	out_data_0,
	Selector6,
	Selector5)/* synthesis synthesis_greybox=0 */;
input 	h2f_WLAST_0;
input 	h2f_ARLEN_0;
input 	h2f_ARLEN_1;
input 	h2f_ARLEN_2;
input 	h2f_ARLEN_3;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWADDR_0;
input 	h2f_AWADDR_1;
input 	h2f_AWADDR_2;
input 	h2f_AWADDR_3;
input 	h2f_AWADDR_4;
input 	h2f_AWADDR_5;
input 	h2f_AWADDR_6;
input 	h2f_AWADDR_7;
input 	h2f_AWADDR_8;
input 	h2f_AWADDR_9;
input 	h2f_AWADDR_10;
input 	h2f_AWADDR_11;
input 	h2f_AWADDR_12;
input 	h2f_AWADDR_13;
input 	h2f_AWADDR_14;
input 	h2f_AWADDR_15;
input 	h2f_AWADDR_16;
input 	h2f_AWADDR_17;
input 	h2f_AWADDR_18;
input 	h2f_AWADDR_19;
input 	h2f_AWADDR_20;
input 	h2f_AWADDR_21;
input 	h2f_AWADDR_22;
input 	h2f_AWADDR_23;
input 	h2f_AWADDR_24;
input 	h2f_AWADDR_25;
input 	h2f_AWADDR_26;
input 	h2f_AWADDR_27;
input 	h2f_AWBURST_0;
input 	h2f_AWBURST_1;
input 	h2f_AWLEN_0;
input 	h2f_AWLEN_1;
input 	h2f_AWLEN_2;
input 	h2f_AWLEN_3;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	outclk_wire_0;
output 	address_burst_24;
output 	address_burst_25;
output 	address_burst_23;
output 	address_burst_13;
output 	address_burst_21;
output 	address_burst_22;
output 	address_burst_19;
output 	address_burst_20;
output 	address_burst_15;
output 	address_burst_16;
output 	address_burst_17;
output 	address_burst_18;
output 	address_burst_26;
output 	address_burst_27;
output 	address_burst_12;
output 	address_burst_14;
output 	address_burst_10;
output 	address_burst_11;
output 	address_burst_9;
output 	address_burst_8;
output 	Add4;
output 	Add5;
output 	Add41;
output 	Add51;
output 	Add42;
output 	Add52;
output 	Add43;
output 	Add53;
output 	Add44;
output 	Add54;
output 	Add55;
output 	Add45;
output 	Add56;
output 	Add46;
output 	Add47;
output 	Add57;
output 	Add48;
output 	Add58;
input 	in_ready;
input 	nxt_in_ready;
output 	sop_enable1;
output 	address_burst_7;
output 	address_burst_6;
output 	address_burst_2;
output 	address_burst_3;
output 	address_burst_4;
output 	address_burst_5;
input 	sink_ready;
input 	sink_ready1;
input 	cmd_sink_ready;
input 	last_cycle;
output 	awready;
input 	last_cycle1;
output 	wready;
output 	LessThan11;
output 	Add3;
output 	log2ceil;
output 	address_burst_1;
output 	LessThan10;
output 	Add31;
output 	address_burst_0;
output 	out_data_2;
output 	out_data_3;
output 	burst_bytecount_4;
output 	burst_bytecount_6;
output 	burst_bytecount_5;
output 	burst_bytecount_7;
output 	Add0;
output 	Add2;
output 	Add01;
output 	Add21;
output 	Add22;
output 	write_cp_data_188;
output 	write_cp_data_187;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_data_7;
output 	Add1;
output 	out_data_9;
output 	out_data_6;
output 	LessThan16;
output 	out_data_8;
output 	LessThan12;
output 	Selector26;
output 	out_data_4;
output 	LessThan14;
output 	out_data_5;
output 	LessThan15;
output 	LessThan2;
output 	Add32;
output 	Selector7;
output 	out_data_1;
output 	Decoder0;
output 	Selector8;
output 	out_data_0;
output 	Selector6;
output 	Selector5;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|Decoder0~0_combout ;
wire \align_address_to_size|Decoder0~2_combout ;
wire \align_address_to_size|Decoder0~3_combout ;
wire \align_address_to_size|Decoder0~4_combout ;
wire \align_address_to_size|Decoder0~5_combout ;
wire \align_address_to_size|Decoder0~6_combout ;
wire \align_address_to_size|Decoder0~7_combout ;
wire \Add4~2 ;
wire \Add5~2 ;
wire \Add4~6 ;
wire \Add5~6 ;
wire \Add4~10 ;
wire \Add5~10 ;
wire \Add4~14 ;
wire \Add5~14 ;
wire \Add4~18 ;
wire \Add5~18 ;
wire \Add5~22 ;
wire \Add4~22 ;
wire \Add5~26 ;
wire \Add4~26 ;
wire \Add4~30 ;
wire \Add5~30 ;
wire \Decoder1~0_combout ;
wire \Decoder1~1_combout ;
wire \Decoder1~2_combout ;
wire \Decoder1~3_combout ;
wire \Decoder1~4_combout ;
wire \Decoder1~5_combout ;
wire \Decoder1~6_combout ;
wire \Decoder1~7_combout ;
wire \sop_enable~0_combout ;
wire \Add1~0_combout ;
wire \Add1~1_combout ;
wire \Add1~2_combout ;
wire \write_cp_data[184]~2_combout ;
wire \write_cp_data[186]~3_combout ;
wire \write_cp_data[185]~4_combout ;
wire \Add7~0_combout ;
wire \Add7~1_combout ;
wire \Add7~2_combout ;
wire \Add7~3_combout ;
wire \burst_bytecount[8]~q ;


Computer_System_altera_merlin_address_alignment align_address_to_size(
	.h2f_AWADDR_0(h2f_AWADDR_0),
	.h2f_AWADDR_1(h2f_AWADDR_1),
	.h2f_AWADDR_2(h2f_AWADDR_2),
	.h2f_AWADDR_3(h2f_AWADDR_3),
	.h2f_AWADDR_4(h2f_AWADDR_4),
	.h2f_AWADDR_5(h2f_AWADDR_5),
	.h2f_AWADDR_6(h2f_AWADDR_6),
	.h2f_AWADDR_7(h2f_AWADDR_7),
	.h2f_AWADDR_8(h2f_AWADDR_8),
	.h2f_AWADDR_9(h2f_AWADDR_9),
	.h2f_AWADDR_10(h2f_AWADDR_10),
	.h2f_AWADDR_11(h2f_AWADDR_11),
	.h2f_AWADDR_12(h2f_AWADDR_12),
	.h2f_AWADDR_13(h2f_AWADDR_13),
	.h2f_AWADDR_14(h2f_AWADDR_14),
	.h2f_AWADDR_15(h2f_AWADDR_15),
	.h2f_AWADDR_16(h2f_AWADDR_16),
	.h2f_AWADDR_17(h2f_AWADDR_17),
	.h2f_AWADDR_18(h2f_AWADDR_18),
	.h2f_AWADDR_19(h2f_AWADDR_19),
	.h2f_AWADDR_20(h2f_AWADDR_20),
	.h2f_AWADDR_21(h2f_AWADDR_21),
	.h2f_AWADDR_22(h2f_AWADDR_22),
	.h2f_AWADDR_23(h2f_AWADDR_23),
	.h2f_AWADDR_24(h2f_AWADDR_24),
	.h2f_AWADDR_25(h2f_AWADDR_25),
	.h2f_AWADDR_26(h2f_AWADDR_26),
	.h2f_AWADDR_27(h2f_AWADDR_27),
	.h2f_AWBURST_0(h2f_AWBURST_0),
	.h2f_AWBURST_1(h2f_AWBURST_1),
	.h2f_AWLEN_3(h2f_AWLEN_3),
	.h2f_AWSIZE_0(h2f_AWSIZE_0),
	.h2f_AWSIZE_1(h2f_AWSIZE_1),
	.h2f_AWSIZE_2(h2f_AWSIZE_2),
	.clk(outclk_wire_0),
	.address_burst_24(address_burst_24),
	.address_burst_25(address_burst_25),
	.address_burst_23(address_burst_23),
	.address_burst_13(address_burst_13),
	.address_burst_21(address_burst_21),
	.address_burst_22(address_burst_22),
	.address_burst_19(address_burst_19),
	.address_burst_20(address_burst_20),
	.address_burst_15(address_burst_15),
	.address_burst_16(address_burst_16),
	.address_burst_17(address_burst_17),
	.address_burst_18(address_burst_18),
	.address_burst_26(address_burst_26),
	.address_burst_27(address_burst_27),
	.address_burst_12(address_burst_12),
	.address_burst_14(address_burst_14),
	.address_burst_10(address_burst_10),
	.address_burst_11(address_burst_11),
	.address_burst_9(address_burst_9),
	.address_burst_8(address_burst_8),
	.sop_enable(sop_enable1),
	.address_burst_7(address_burst_7),
	.address_burst_6(address_burst_6),
	.address_burst_2(address_burst_2),
	.address_burst_3(address_burst_3),
	.address_burst_4(address_burst_4),
	.address_burst_5(address_burst_5),
	.wready(wready),
	.Add1(\Add1~0_combout ),
	.LessThan11(LessThan11),
	.address_burst_1(address_burst_1),
	.LessThan10(LessThan10),
	.address_burst_0(address_burst_0),
	.out_data_2(out_data_2),
	.out_data_3(out_data_3),
	.reset(altera_reset_synchronizer_int_chain_out),
	.out_data_7(out_data_7),
	.Add11(Add1),
	.out_data_9(out_data_9),
	.out_data_6(out_data_6),
	.LessThan16(LessThan16),
	.out_data_8(out_data_8),
	.LessThan12(LessThan12),
	.Selector26(Selector26),
	.out_data_4(out_data_4),
	.LessThan14(LessThan14),
	.out_data_5(out_data_5),
	.LessThan15(LessThan15),
	.LessThan2(LessThan2),
	.Decoder0(\align_address_to_size|Decoder0~0_combout ),
	.out_data_1(out_data_1),
	.Decoder01(Decoder0),
	.out_data_0(out_data_0),
	.Decoder02(\align_address_to_size|Decoder0~2_combout ),
	.Decoder03(\align_address_to_size|Decoder0~3_combout ),
	.Decoder04(\align_address_to_size|Decoder0~4_combout ),
	.Decoder05(\align_address_to_size|Decoder0~5_combout ),
	.Decoder06(\align_address_to_size|Decoder0~6_combout ),
	.Decoder07(\align_address_to_size|Decoder0~7_combout ));

cyclonev_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add4),
	.cout(\Add4~2 ),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h00000000000000FF;
defparam \Add4~1 .shared_arith = "off";

cyclonev_lcell_comb \Add5~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add5),
	.cout(\Add5~2 ),
	.shareout());
defparam \Add5~1 .extended_lut = "off";
defparam \Add5~1 .lut_mask = 64'h00000000000000FF;
defparam \Add5~1 .shared_arith = "off";

cyclonev_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add41),
	.cout(\Add4~6 ),
	.shareout());
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h00000000000000FF;
defparam \Add4~5 .shared_arith = "off";

cyclonev_lcell_comb \Add5~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add51),
	.cout(\Add5~6 ),
	.shareout());
defparam \Add5~5 .extended_lut = "off";
defparam \Add5~5 .lut_mask = 64'h00000000000000FF;
defparam \Add5~5 .shared_arith = "off";

cyclonev_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add42),
	.cout(\Add4~10 ),
	.shareout());
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h00000000000000FF;
defparam \Add4~9 .shared_arith = "off";

cyclonev_lcell_comb \Add5~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add52),
	.cout(\Add5~10 ),
	.shareout());
defparam \Add5~9 .extended_lut = "off";
defparam \Add5~9 .lut_mask = 64'h00000000000000FF;
defparam \Add5~9 .shared_arith = "off";

cyclonev_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add43),
	.cout(\Add4~14 ),
	.shareout());
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h00000000000000FF;
defparam \Add4~13 .shared_arith = "off";

cyclonev_lcell_comb \Add5~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add53),
	.cout(\Add5~14 ),
	.shareout());
defparam \Add5~13 .extended_lut = "off";
defparam \Add5~13 .lut_mask = 64'h00000000000000FF;
defparam \Add5~13 .shared_arith = "off";

cyclonev_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add44),
	.cout(\Add4~18 ),
	.shareout());
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h00000000000000FF;
defparam \Add4~17 .shared_arith = "off";

cyclonev_lcell_comb \Add5~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add54),
	.cout(\Add5~18 ),
	.shareout());
defparam \Add5~17 .extended_lut = "off";
defparam \Add5~17 .lut_mask = 64'h00000000000000FF;
defparam \Add5~17 .shared_arith = "off";

cyclonev_lcell_comb \Add5~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add55),
	.cout(\Add5~22 ),
	.shareout());
defparam \Add5~21 .extended_lut = "off";
defparam \Add5~21 .lut_mask = 64'h00000000000000FF;
defparam \Add5~21 .shared_arith = "off";

cyclonev_lcell_comb \Add4~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add45),
	.cout(\Add4~22 ),
	.shareout());
defparam \Add4~21 .extended_lut = "off";
defparam \Add4~21 .lut_mask = 64'h00000000000000FF;
defparam \Add4~21 .shared_arith = "off";

cyclonev_lcell_comb \Add5~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add56),
	.cout(\Add5~26 ),
	.shareout());
defparam \Add5~25 .extended_lut = "off";
defparam \Add5~25 .lut_mask = 64'h00000000000000FF;
defparam \Add5~25 .shared_arith = "off";

cyclonev_lcell_comb \Add4~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add46),
	.cout(\Add4~26 ),
	.shareout());
defparam \Add4~25 .extended_lut = "off";
defparam \Add4~25 .lut_mask = 64'h00000000000000FF;
defparam \Add4~25 .shared_arith = "off";

cyclonev_lcell_comb \Add4~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add47),
	.cout(\Add4~30 ),
	.shareout());
defparam \Add4~29 .extended_lut = "off";
defparam \Add4~29 .lut_mask = 64'h00000000000000FF;
defparam \Add4~29 .shared_arith = "off";

cyclonev_lcell_comb \Add5~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add57),
	.cout(\Add5~30 ),
	.shareout());
defparam \Add5~29 .extended_lut = "off";
defparam \Add5~29 .lut_mask = 64'h00000000000000FF;
defparam \Add5~29 .shared_arith = "off";

cyclonev_lcell_comb \Add4~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add48),
	.cout(),
	.shareout());
defparam \Add4~33 .extended_lut = "off";
defparam \Add4~33 .lut_mask = 64'h0000FFFF0000FFFF;
defparam \Add4~33 .shared_arith = "off";

cyclonev_lcell_comb \Add5~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add58),
	.cout(),
	.shareout());
defparam \Add5~33 .extended_lut = "off";
defparam \Add5~33 .lut_mask = 64'h0000FFFF0000FFFF;
defparam \Add5~33 .shared_arith = "off";

dffeas sop_enable(
	.clk(outclk_wire_0),
	.d(\sop_enable~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(sop_enable1),
	.prn(vcc));
defparam sop_enable.is_wysiwyg = "true";
defparam sop_enable.power_up = "low";

cyclonev_lcell_comb \awready~0 (
	.dataa(!in_ready),
	.datab(!nxt_in_ready),
	.datac(!sink_ready),
	.datad(!sink_ready1),
	.datae(!cmd_sink_ready),
	.dataf(!last_cycle),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(awready),
	.sumout(),
	.cout(),
	.shareout());
defparam \awready~0 .extended_lut = "off";
defparam \awready~0 .lut_mask = 64'h0000000008FF0000;
defparam \awready~0 .shared_arith = "off";

cyclonev_lcell_comb \wready~0 (
	.dataa(!in_ready),
	.datab(!nxt_in_ready),
	.datac(!sink_ready),
	.datad(!sink_ready1),
	.datae(!cmd_sink_ready),
	.dataf(!last_cycle1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wready),
	.sumout(),
	.cout(),
	.shareout());
defparam \wready~0 .extended_lut = "off";
defparam \wready~0 .lut_mask = 64'h0000000008FF0000;
defparam \wready~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan11~0 (
	.dataa(!h2f_AWLEN_3),
	.datab(!h2f_AWSIZE_2),
	.datac(!\Add1~0_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan11),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan11~0 .extended_lut = "off";
defparam \LessThan11~0 .lut_mask = 64'h8000800080008000;
defparam \LessThan11~0 .shared_arith = "off";

cyclonev_lcell_comb \Add3~0 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!h2f_ARLEN_3),
	.datae(!h2f_ARSIZE_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~0 .extended_lut = "off";
defparam \Add3~0 .lut_mask = 64'h00004F0000004F00;
defparam \Add3~0 .shared_arith = "off";

cyclonev_lcell_comb \log2ceil~0 (
	.dataa(!h2f_ARLEN_1),
	.datab(!h2f_ARLEN_2),
	.datac(!h2f_ARLEN_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(log2ceil),
	.sumout(),
	.cout(),
	.shareout());
defparam \log2ceil~0 .extended_lut = "off";
defparam \log2ceil~0 .lut_mask = 64'h7070707070707070;
defparam \log2ceil~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan10~0 (
	.dataa(!h2f_AWLEN_3),
	.datab(!h2f_AWSIZE_2),
	.datac(!\Add1~0_combout ),
	.datad(!\Add1~1_combout ),
	.datae(!\Add1~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan10),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan10~0 .extended_lut = "off";
defparam \LessThan10~0 .lut_mask = 64'h8000000080000000;
defparam \LessThan10~0 .shared_arith = "off";

cyclonev_lcell_comb \Add3~1 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!h2f_ARLEN_3),
	.datae(!h2f_ARSIZE_0),
	.dataf(!h2f_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add31),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h00000F003F007F00;
defparam \Add3~1 .shared_arith = "off";

dffeas \burst_bytecount[4] (
	.clk(outclk_wire_0),
	.d(\write_cp_data[184]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_4),
	.prn(vcc));
defparam \burst_bytecount[4] .is_wysiwyg = "true";
defparam \burst_bytecount[4] .power_up = "low";

dffeas \burst_bytecount[6] (
	.clk(outclk_wire_0),
	.d(\Add7~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_6),
	.prn(vcc));
defparam \burst_bytecount[6] .is_wysiwyg = "true";
defparam \burst_bytecount[6] .power_up = "low";

dffeas \burst_bytecount[5] (
	.clk(outclk_wire_0),
	.d(\Add7~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_5),
	.prn(vcc));
defparam \burst_bytecount[5] .is_wysiwyg = "true";
defparam \burst_bytecount[5] .power_up = "low";

dffeas \burst_bytecount[7] (
	.clk(outclk_wire_0),
	.d(\Add7~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_7),
	.prn(vcc));
defparam \burst_bytecount[7] .is_wysiwyg = "true";
defparam \burst_bytecount[7] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!h2f_AWLEN_2),
	.datad(!h2f_AWLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h01FE01FE01FE01FE;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add2~0 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!h2f_ARLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~0 .extended_lut = "off";
defparam \Add2~0 .lut_mask = 64'h01FE01FE01FE01FE;
defparam \Add2~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!h2f_AWLEN_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add01),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h1E1E1E1E1E1E1E1E;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add21),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h1E1E1E1E1E1E1E1E;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \Add2~2 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add22),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~2 .extended_lut = "off";
defparam \Add2~2 .lut_mask = 64'h6666666666666666;
defparam \Add2~2 .shared_arith = "off";

cyclonev_lcell_comb \write_cp_data[188]~0 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!h2f_AWLEN_2),
	.datad(!h2f_AWLEN_3),
	.datae(!sop_enable1),
	.dataf(!\burst_bytecount[8]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_188),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[188]~0 .extended_lut = "off";
defparam \write_cp_data[188]~0 .lut_mask = 64'h000100000001FFFF;
defparam \write_cp_data[188]~0 .shared_arith = "off";

cyclonev_lcell_comb \write_cp_data[187]~1 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!h2f_AWLEN_2),
	.datad(!h2f_AWLEN_3),
	.datae(!sop_enable1),
	.dataf(!burst_bytecount_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_187),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[187]~1 .extended_lut = "off";
defparam \write_cp_data[187]~1 .lut_mask = 64'h01FE000001FEFFFF;
defparam \write_cp_data[187]~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~3 (
	.dataa(!h2f_AWLEN_3),
	.datab(!h2f_AWSIZE_2),
	.datac(!\Add1~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~3 .extended_lut = "off";
defparam \Add1~3 .lut_mask = 64'h1717171717171717;
defparam \Add1~3 .shared_arith = "off";

cyclonev_lcell_comb \LessThan16~0 (
	.dataa(!h2f_AWLEN_3),
	.datab(!h2f_AWSIZE_2),
	.datac(!\Add1~0_combout ),
	.datad(!\Add1~1_combout ),
	.datae(!\Add1~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan16),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan16~0 .extended_lut = "off";
defparam \LessThan16~0 .lut_mask = 64'hE8E8E880E8E8E880;
defparam \LessThan16~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan12~0 (
	.dataa(!h2f_AWLEN_3),
	.datab(!h2f_AWSIZE_2),
	.datac(!\Add1~0_combout ),
	.datad(!\Add1~1_combout ),
	.datae(!\Add1~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan12),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan12~0 .extended_lut = "off";
defparam \LessThan12~0 .lut_mask = 64'h8080800080808000;
defparam \LessThan12~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan14~0 (
	.dataa(!h2f_AWLEN_3),
	.datab(!h2f_AWSIZE_2),
	.datac(!\Add1~0_combout ),
	.datad(!\Add1~1_combout ),
	.datae(!\Add1~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan14),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan14~0 .extended_lut = "off";
defparam \LessThan14~0 .lut_mask = 64'hE8808080E8808080;
defparam \LessThan14~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan15~0 (
	.dataa(!h2f_AWLEN_3),
	.datab(!h2f_AWSIZE_2),
	.datac(!\Add1~0_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan15),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan15~0 .extended_lut = "off";
defparam \LessThan15~0 .lut_mask = 64'hE880E880E880E880;
defparam \LessThan15~0 .shared_arith = "off";

cyclonev_lcell_comb \Add3~2 (
	.dataa(!h2f_ARLEN_3),
	.datab(!h2f_ARSIZE_2),
	.datac(!Add31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add32),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~2 .extended_lut = "off";
defparam \Add3~2 .lut_mask = 64'h1717171717171717;
defparam \Add3~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector7~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!LessThan11),
	.datad(!Add4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector7),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'h8A028A028A028A02;
defparam \Selector7~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!LessThan10),
	.datad(!Add41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector8),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'h8A028A028A028A02;
defparam \Selector8~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!LessThan12),
	.datad(!Add42),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector6),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'h8A028A028A028A02;
defparam \Selector6~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!Add43),
	.datad(!h2f_AWLEN_3),
	.datae(!h2f_AWSIZE_2),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector5),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'hA280808080808080;
defparam \Selector5~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~0 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~0 .extended_lut = "off";
defparam \Decoder1~0 .lut_mask = 64'h4040404040404040;
defparam \Decoder1~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~1 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~1 .extended_lut = "off";
defparam \Decoder1~1 .lut_mask = 64'h8080808080808080;
defparam \Decoder1~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~2 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~2 .extended_lut = "off";
defparam \Decoder1~2 .lut_mask = 64'h2020202020202020;
defparam \Decoder1~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~3 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~3 .extended_lut = "off";
defparam \Decoder1~3 .lut_mask = 64'h1010101010101010;
defparam \Decoder1~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~4 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~4 .extended_lut = "off";
defparam \Decoder1~4 .lut_mask = 64'h0808080808080808;
defparam \Decoder1~4 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~5 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~5 .extended_lut = "off";
defparam \Decoder1~5 .lut_mask = 64'h0404040404040404;
defparam \Decoder1~5 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~6 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~6 .extended_lut = "off";
defparam \Decoder1~6 .lut_mask = 64'h0202020202020202;
defparam \Decoder1~6 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~7 (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~7 .extended_lut = "off";
defparam \Decoder1~7 .lut_mask = 64'h0101010101010101;
defparam \Decoder1~7 .shared_arith = "off";

cyclonev_lcell_comb \sop_enable~0 (
	.dataa(!h2f_WLAST_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sop_enable~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sop_enable~0 .extended_lut = "off";
defparam \sop_enable~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sop_enable~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!h2f_AWLEN_2),
	.datad(!h2f_AWLEN_3),
	.datae(!h2f_AWSIZE_0),
	.dataf(!h2f_AWSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h00000F003F007F00;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!h2f_AWLEN_2),
	.datad(!h2f_AWLEN_3),
	.datae(!h2f_AWSIZE_0),
	.dataf(!h2f_AWSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h3F007000C0FF8FFF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~2 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!h2f_AWLEN_2),
	.datad(!h2f_AWLEN_3),
	.datae(!h2f_AWSIZE_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~2 .extended_lut = "off";
defparam \Add1~2 .lut_mask = 64'h4F00B0FF4F00B0FF;
defparam \Add1~2 .shared_arith = "off";

cyclonev_lcell_comb \write_cp_data[184]~2 (
	.dataa(!h2f_AWLEN_0),
	.datab(!sop_enable1),
	.datac(!burst_bytecount_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_cp_data[184]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[184]~2 .extended_lut = "off";
defparam \write_cp_data[184]~2 .lut_mask = 64'h7474747474747474;
defparam \write_cp_data[184]~2 .shared_arith = "off";

cyclonev_lcell_comb \write_cp_data[186]~3 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!h2f_AWLEN_2),
	.datad(!sop_enable1),
	.datae(!burst_bytecount_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_cp_data[186]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[186]~3 .extended_lut = "off";
defparam \write_cp_data[186]~3 .lut_mask = 64'h1E001EFF1E001EFF;
defparam \write_cp_data[186]~3 .shared_arith = "off";

cyclonev_lcell_comb \write_cp_data[185]~4 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!sop_enable1),
	.datad(!burst_bytecount_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_cp_data[185]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[185]~4 .extended_lut = "off";
defparam \write_cp_data[185]~4 .lut_mask = 64'h606F606F606F606F;
defparam \write_cp_data[185]~4 .shared_arith = "off";

cyclonev_lcell_comb \Add7~0 (
	.dataa(!\write_cp_data[184]~2_combout ),
	.datab(!\write_cp_data[186]~3_combout ),
	.datac(!\write_cp_data[185]~4_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~0 .extended_lut = "off";
defparam \Add7~0 .lut_mask = 64'h6363636363636363;
defparam \Add7~0 .shared_arith = "off";

cyclonev_lcell_comb \Add7~1 (
	.dataa(!\write_cp_data[184]~2_combout ),
	.datab(!\write_cp_data[185]~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h6666666666666666;
defparam \Add7~1 .shared_arith = "off";

cyclonev_lcell_comb \Add7~2 (
	.dataa(!\write_cp_data[184]~2_combout ),
	.datab(!\write_cp_data[186]~3_combout ),
	.datac(!\write_cp_data[185]~4_combout ),
	.datad(!write_cp_data_187),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~2 .extended_lut = "off";
defparam \Add7~2 .lut_mask = 64'h40BF40BF40BF40BF;
defparam \Add7~2 .shared_arith = "off";

cyclonev_lcell_comb \Add7~3 (
	.dataa(!\write_cp_data[184]~2_combout ),
	.datab(!\write_cp_data[186]~3_combout ),
	.datac(!\write_cp_data[185]~4_combout ),
	.datad(!write_cp_data_187),
	.datae(!write_cp_data_188),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~3 .extended_lut = "off";
defparam \Add7~3 .lut_mask = 64'h4000BFFF4000BFFF;
defparam \Add7~3 .shared_arith = "off";

dffeas \burst_bytecount[8] (
	.clk(outclk_wire_0),
	.d(\Add7~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\burst_bytecount[8]~q ),
	.prn(vcc));
defparam \burst_bytecount[8] .is_wysiwyg = "true";
defparam \burst_bytecount[8] .power_up = "low";

endmodule

module Computer_System_altera_merlin_address_alignment (
	h2f_AWADDR_0,
	h2f_AWADDR_1,
	h2f_AWADDR_2,
	h2f_AWADDR_3,
	h2f_AWADDR_4,
	h2f_AWADDR_5,
	h2f_AWADDR_6,
	h2f_AWADDR_7,
	h2f_AWADDR_8,
	h2f_AWADDR_9,
	h2f_AWADDR_10,
	h2f_AWADDR_11,
	h2f_AWADDR_12,
	h2f_AWADDR_13,
	h2f_AWADDR_14,
	h2f_AWADDR_15,
	h2f_AWADDR_16,
	h2f_AWADDR_17,
	h2f_AWADDR_18,
	h2f_AWADDR_19,
	h2f_AWADDR_20,
	h2f_AWADDR_21,
	h2f_AWADDR_22,
	h2f_AWADDR_23,
	h2f_AWADDR_24,
	h2f_AWADDR_25,
	h2f_AWADDR_26,
	h2f_AWADDR_27,
	h2f_AWBURST_0,
	h2f_AWBURST_1,
	h2f_AWLEN_3,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	clk,
	address_burst_24,
	address_burst_25,
	address_burst_23,
	address_burst_13,
	address_burst_21,
	address_burst_22,
	address_burst_19,
	address_burst_20,
	address_burst_15,
	address_burst_16,
	address_burst_17,
	address_burst_18,
	address_burst_26,
	address_burst_27,
	address_burst_12,
	address_burst_14,
	address_burst_10,
	address_burst_11,
	address_burst_9,
	address_burst_8,
	sop_enable,
	address_burst_7,
	address_burst_6,
	address_burst_2,
	address_burst_3,
	address_burst_4,
	address_burst_5,
	wready,
	Add1,
	LessThan11,
	address_burst_1,
	LessThan10,
	address_burst_0,
	out_data_2,
	out_data_3,
	reset,
	out_data_7,
	Add11,
	out_data_9,
	out_data_6,
	LessThan16,
	out_data_8,
	LessThan12,
	Selector26,
	out_data_4,
	LessThan14,
	out_data_5,
	LessThan15,
	LessThan2,
	Decoder0,
	out_data_1,
	Decoder01,
	out_data_0,
	Decoder02,
	Decoder03,
	Decoder04,
	Decoder05,
	Decoder06,
	Decoder07)/* synthesis synthesis_greybox=0 */;
input 	h2f_AWADDR_0;
input 	h2f_AWADDR_1;
input 	h2f_AWADDR_2;
input 	h2f_AWADDR_3;
input 	h2f_AWADDR_4;
input 	h2f_AWADDR_5;
input 	h2f_AWADDR_6;
input 	h2f_AWADDR_7;
input 	h2f_AWADDR_8;
input 	h2f_AWADDR_9;
input 	h2f_AWADDR_10;
input 	h2f_AWADDR_11;
input 	h2f_AWADDR_12;
input 	h2f_AWADDR_13;
input 	h2f_AWADDR_14;
input 	h2f_AWADDR_15;
input 	h2f_AWADDR_16;
input 	h2f_AWADDR_17;
input 	h2f_AWADDR_18;
input 	h2f_AWADDR_19;
input 	h2f_AWADDR_20;
input 	h2f_AWADDR_21;
input 	h2f_AWADDR_22;
input 	h2f_AWADDR_23;
input 	h2f_AWADDR_24;
input 	h2f_AWADDR_25;
input 	h2f_AWADDR_26;
input 	h2f_AWADDR_27;
input 	h2f_AWBURST_0;
input 	h2f_AWBURST_1;
input 	h2f_AWLEN_3;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	clk;
output 	address_burst_24;
output 	address_burst_25;
output 	address_burst_23;
output 	address_burst_13;
output 	address_burst_21;
output 	address_burst_22;
output 	address_burst_19;
output 	address_burst_20;
output 	address_burst_15;
output 	address_burst_16;
output 	address_burst_17;
output 	address_burst_18;
output 	address_burst_26;
output 	address_burst_27;
output 	address_burst_12;
output 	address_burst_14;
output 	address_burst_10;
output 	address_burst_11;
output 	address_burst_9;
output 	address_burst_8;
input 	sop_enable;
output 	address_burst_7;
output 	address_burst_6;
output 	address_burst_2;
output 	address_burst_3;
output 	address_burst_4;
output 	address_burst_5;
input 	wready;
input 	Add1;
input 	LessThan11;
output 	address_burst_1;
input 	LessThan10;
output 	address_burst_0;
output 	out_data_2;
output 	out_data_3;
input 	reset;
output 	out_data_7;
input 	Add11;
output 	out_data_9;
output 	out_data_6;
input 	LessThan16;
output 	out_data_8;
input 	LessThan12;
output 	Selector26;
output 	out_data_4;
input 	LessThan14;
output 	out_data_5;
input 	LessThan15;
output 	LessThan2;
output 	Decoder0;
output 	out_data_1;
output 	Decoder01;
output 	out_data_0;
output 	Decoder02;
output 	Decoder03;
output 	Decoder04;
output 	Decoder05;
output 	Decoder06;
output 	Decoder07;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \aligned_address_bits[3]~combout ;
wire \aligned_address_bits[1]~combout ;
wire \Add0~110 ;
wire \Add0~106 ;
wire \Add0~90 ;
wire \Add0~94 ;
wire \Add0~98 ;
wire \Add0~102 ;
wire \Add0~82 ;
wire \Add0~74 ;
wire \Add0~86 ;
wire \Add0~78 ;
wire \Add0~66 ;
wire \Add0~70 ;
wire \Add0~58 ;
wire \Add0~14 ;
wire \Add0~62 ;
wire \Add0~34 ;
wire \Add0~38 ;
wire \Add0~42 ;
wire \Add0~46 ;
wire \Add0~26 ;
wire \Add0~30 ;
wire \Add0~18 ;
wire \Add0~22 ;
wire \Add0~10 ;
wire \Add0~1_sumout ;
wire \out_data[24]~2_combout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \out_data[25]~3_combout ;
wire \Add0~9_sumout ;
wire \out_data[23]~4_combout ;
wire \Add0~13_sumout ;
wire \out_data[13]~5_combout ;
wire \Add0~17_sumout ;
wire \out_data[21]~6_combout ;
wire \Add0~21_sumout ;
wire \out_data[22]~7_combout ;
wire \Add0~25_sumout ;
wire \out_data[19]~8_combout ;
wire \Add0~29_sumout ;
wire \out_data[20]~9_combout ;
wire \Add0~33_sumout ;
wire \out_data[15]~10_combout ;
wire \Add0~37_sumout ;
wire \out_data[16]~11_combout ;
wire \Add0~41_sumout ;
wire \out_data[17]~12_combout ;
wire \Add0~45_sumout ;
wire \out_data[18]~13_combout ;
wire \Add0~6 ;
wire \Add0~49_sumout ;
wire \out_data[26]~14_combout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \out_data[27]~15_combout ;
wire \Add0~57_sumout ;
wire \out_data[12]~16_combout ;
wire \Add0~61_sumout ;
wire \out_data[14]~17_combout ;
wire \Add0~65_sumout ;
wire \out_data[10]~18_combout ;
wire \Add0~69_sumout ;
wire \out_data[11]~19_combout ;
wire \Add0~77_sumout ;
wire \Add0~85_sumout ;
wire \Add1~30 ;
wire \Add1~26 ;
wire \Add1~10 ;
wire \Add1~14 ;
wire \Add1~18 ;
wire \Add1~22 ;
wire \Add1~6 ;
wire \Add1~1_sumout ;
wire \Add0~73_sumout ;
wire \Selector22~0_combout ;
wire \Add1~5_sumout ;
wire \Add0~81_sumout ;
wire \Selector23~0_combout ;
wire \Add1~9_sumout ;
wire \Add0~89_sumout ;
wire \Selector27~0_combout ;
wire \Add1~13_sumout ;
wire \Add0~93_sumout ;
wire \Selector26~1_combout ;
wire \Add1~17_sumout ;
wire \Add0~97_sumout ;
wire \Selector25~0_combout ;
wire \Add1~21_sumout ;
wire \Add0~101_sumout ;
wire \Selector24~0_combout ;
wire \Add1~25_sumout ;
wire \Add0~105_sumout ;
wire \Selector28~0_combout ;
wire \Add1~29_sumout ;
wire \Add0~109_sumout ;
wire \Selector29~0_combout ;


dffeas \address_burst[24] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(\out_data[24]~2_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_24),
	.prn(vcc));
defparam \address_burst[24] .is_wysiwyg = "true";
defparam \address_burst[24] .power_up = "low";

dffeas \address_burst[25] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(\out_data[25]~3_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_25),
	.prn(vcc));
defparam \address_burst[25] .is_wysiwyg = "true";
defparam \address_burst[25] .power_up = "low";

dffeas \address_burst[23] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(\out_data[23]~4_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_23),
	.prn(vcc));
defparam \address_burst[23] .is_wysiwyg = "true";
defparam \address_burst[23] .power_up = "low";

dffeas \address_burst[13] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(\out_data[13]~5_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_13),
	.prn(vcc));
defparam \address_burst[13] .is_wysiwyg = "true";
defparam \address_burst[13] .power_up = "low";

dffeas \address_burst[21] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(\out_data[21]~6_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_21),
	.prn(vcc));
defparam \address_burst[21] .is_wysiwyg = "true";
defparam \address_burst[21] .power_up = "low";

dffeas \address_burst[22] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(\out_data[22]~7_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_22),
	.prn(vcc));
defparam \address_burst[22] .is_wysiwyg = "true";
defparam \address_burst[22] .power_up = "low";

dffeas \address_burst[19] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(\out_data[19]~8_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_19),
	.prn(vcc));
defparam \address_burst[19] .is_wysiwyg = "true";
defparam \address_burst[19] .power_up = "low";

dffeas \address_burst[20] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(\out_data[20]~9_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_20),
	.prn(vcc));
defparam \address_burst[20] .is_wysiwyg = "true";
defparam \address_burst[20] .power_up = "low";

dffeas \address_burst[15] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(\out_data[15]~10_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_15),
	.prn(vcc));
defparam \address_burst[15] .is_wysiwyg = "true";
defparam \address_burst[15] .power_up = "low";

dffeas \address_burst[16] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(\out_data[16]~11_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_16),
	.prn(vcc));
defparam \address_burst[16] .is_wysiwyg = "true";
defparam \address_burst[16] .power_up = "low";

dffeas \address_burst[17] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(\out_data[17]~12_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_17),
	.prn(vcc));
defparam \address_burst[17] .is_wysiwyg = "true";
defparam \address_burst[17] .power_up = "low";

dffeas \address_burst[18] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(\out_data[18]~13_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_18),
	.prn(vcc));
defparam \address_burst[18] .is_wysiwyg = "true";
defparam \address_burst[18] .power_up = "low";

dffeas \address_burst[26] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(\out_data[26]~14_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_26),
	.prn(vcc));
defparam \address_burst[26] .is_wysiwyg = "true";
defparam \address_burst[26] .power_up = "low";

dffeas \address_burst[27] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(\out_data[27]~15_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_27),
	.prn(vcc));
defparam \address_burst[27] .is_wysiwyg = "true";
defparam \address_burst[27] .power_up = "low";

dffeas \address_burst[12] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(\out_data[12]~16_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_12),
	.prn(vcc));
defparam \address_burst[12] .is_wysiwyg = "true";
defparam \address_burst[12] .power_up = "low";

dffeas \address_burst[14] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(\out_data[14]~17_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_14),
	.prn(vcc));
defparam \address_burst[14] .is_wysiwyg = "true";
defparam \address_burst[14] .power_up = "low";

dffeas \address_burst[10] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(\out_data[10]~18_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_10),
	.prn(vcc));
defparam \address_burst[10] .is_wysiwyg = "true";
defparam \address_burst[10] .power_up = "low";

dffeas \address_burst[11] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(\out_data[11]~19_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_11),
	.prn(vcc));
defparam \address_burst[11] .is_wysiwyg = "true";
defparam \address_burst[11] .power_up = "low";

dffeas \address_burst[9] (
	.clk(clk),
	.d(\Add0~77_sumout ),
	.asdata(out_data_9),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_9),
	.prn(vcc));
defparam \address_burst[9] .is_wysiwyg = "true";
defparam \address_burst[9] .power_up = "low";

dffeas \address_burst[8] (
	.clk(clk),
	.d(\Add0~85_sumout ),
	.asdata(out_data_8),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_AWBURST_0),
	.ena(wready),
	.q(address_burst_8),
	.prn(vcc));
defparam \address_burst[8] .is_wysiwyg = "true";
defparam \address_burst[8] .power_up = "low";

dffeas \address_burst[7] (
	.clk(clk),
	.d(\Selector22~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(address_burst_7),
	.prn(vcc));
defparam \address_burst[7] .is_wysiwyg = "true";
defparam \address_burst[7] .power_up = "low";

dffeas \address_burst[6] (
	.clk(clk),
	.d(\Selector23~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(address_burst_6),
	.prn(vcc));
defparam \address_burst[6] .is_wysiwyg = "true";
defparam \address_burst[6] .power_up = "low";

dffeas \address_burst[2] (
	.clk(clk),
	.d(\Selector27~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(address_burst_2),
	.prn(vcc));
defparam \address_burst[2] .is_wysiwyg = "true";
defparam \address_burst[2] .power_up = "low";

dffeas \address_burst[3] (
	.clk(clk),
	.d(\Selector26~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(address_burst_3),
	.prn(vcc));
defparam \address_burst[3] .is_wysiwyg = "true";
defparam \address_burst[3] .power_up = "low";

dffeas \address_burst[4] (
	.clk(clk),
	.d(\Selector25~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(address_burst_4),
	.prn(vcc));
defparam \address_burst[4] .is_wysiwyg = "true";
defparam \address_burst[4] .power_up = "low";

dffeas \address_burst[5] (
	.clk(clk),
	.d(\Selector24~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(address_burst_5),
	.prn(vcc));
defparam \address_burst[5] .is_wysiwyg = "true";
defparam \address_burst[5] .power_up = "low";

dffeas \address_burst[1] (
	.clk(clk),
	.d(\Selector28~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(address_burst_1),
	.prn(vcc));
defparam \address_burst[1] .is_wysiwyg = "true";
defparam \address_burst[1] .power_up = "low";

dffeas \address_burst[0] (
	.clk(clk),
	.d(\Selector29~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(address_burst_0),
	.prn(vcc));
defparam \address_burst[0] .is_wysiwyg = "true";
defparam \address_burst[0] .power_up = "low";

cyclonev_lcell_comb \out_data[2]~0 (
	.dataa(!h2f_AWADDR_2),
	.datab(!sop_enable),
	.datac(!address_burst_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[2]~0 .extended_lut = "off";
defparam \out_data[2]~0 .lut_mask = 64'h4747474747474747;
defparam \out_data[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[3]~1 (
	.dataa(!h2f_AWADDR_3),
	.datab(!sop_enable),
	.datac(!address_burst_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[3]~1 .extended_lut = "off";
defparam \out_data[3]~1 .lut_mask = 64'h4747474747474747;
defparam \out_data[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[7]~20 (
	.dataa(!h2f_AWADDR_7),
	.datab(!sop_enable),
	.datac(!address_burst_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[7]~20 .extended_lut = "off";
defparam \out_data[7]~20 .lut_mask = 64'h4747474747474747;
defparam \out_data[7]~20 .shared_arith = "off";

cyclonev_lcell_comb \out_data[9]~21 (
	.dataa(!h2f_AWADDR_9),
	.datab(!sop_enable),
	.datac(!address_burst_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[9]~21 .extended_lut = "off";
defparam \out_data[9]~21 .lut_mask = 64'h4747474747474747;
defparam \out_data[9]~21 .shared_arith = "off";

cyclonev_lcell_comb \out_data[6]~22 (
	.dataa(!h2f_AWADDR_6),
	.datab(!sop_enable),
	.datac(!address_burst_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[6]~22 .extended_lut = "off";
defparam \out_data[6]~22 .lut_mask = 64'h4747474747474747;
defparam \out_data[6]~22 .shared_arith = "off";

cyclonev_lcell_comb \out_data[8]~23 (
	.dataa(!h2f_AWADDR_8),
	.datab(!sop_enable),
	.datac(!address_burst_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[8]~23 .extended_lut = "off";
defparam \out_data[8]~23 .lut_mask = 64'h4747474747474747;
defparam \out_data[8]~23 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~0 (
	.dataa(!h2f_AWLEN_3),
	.datab(!h2f_AWSIZE_2),
	.datac(!Add1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector26),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~0 .extended_lut = "off";
defparam \Selector26~0 .lut_mask = 64'h8080808080808080;
defparam \Selector26~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[4]~24 (
	.dataa(!h2f_AWADDR_4),
	.datab(!sop_enable),
	.datac(!address_burst_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[4]~24 .extended_lut = "off";
defparam \out_data[4]~24 .lut_mask = 64'h4747474747474747;
defparam \out_data[4]~24 .shared_arith = "off";

cyclonev_lcell_comb \out_data[5]~25 (
	.dataa(!h2f_AWADDR_5),
	.datab(!sop_enable),
	.datac(!address_burst_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[5]~25 .extended_lut = "off";
defparam \out_data[5]~25 .lut_mask = 64'h4747474747474747;
defparam \out_data[5]~25 .shared_arith = "off";

cyclonev_lcell_comb \LessThan2~0 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan2),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~0 .extended_lut = "off";
defparam \LessThan2~0 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \LessThan2~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'h4040404040404040;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[1]~26 (
	.dataa(!h2f_AWADDR_1),
	.datab(!sop_enable),
	.datac(!address_burst_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[1]~26 .extended_lut = "off";
defparam \out_data[1]~26 .lut_mask = 64'h4747474747474747;
defparam \out_data[1]~26 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder01),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'h8080808080808080;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[0]~27 (
	.dataa(!h2f_AWADDR_0),
	.datab(!sop_enable),
	.datac(!address_burst_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[0]~27 .extended_lut = "off";
defparam \out_data[0]~27 .lut_mask = 64'h4747474747474747;
defparam \out_data[0]~27 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~2 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder02),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~2 .extended_lut = "off";
defparam \Decoder0~2 .lut_mask = 64'h0101010101010101;
defparam \Decoder0~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~3 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder03),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~3 .extended_lut = "off";
defparam \Decoder0~3 .lut_mask = 64'h0202020202020202;
defparam \Decoder0~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~4 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder04),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~4 .extended_lut = "off";
defparam \Decoder0~4 .lut_mask = 64'h2020202020202020;
defparam \Decoder0~4 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~5 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder05),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~5 .extended_lut = "off";
defparam \Decoder0~5 .lut_mask = 64'h1010101010101010;
defparam \Decoder0~5 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~6 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder06),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~6 .extended_lut = "off";
defparam \Decoder0~6 .lut_mask = 64'h0808080808080808;
defparam \Decoder0~6 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~7 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder07),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~7 .extended_lut = "off";
defparam \Decoder0~7 .lut_mask = 64'h0404040404040404;
defparam \Decoder0~7 .shared_arith = "off";

cyclonev_lcell_comb \aligned_address_bits[3] (
	.dataa(!h2f_AWADDR_3),
	.datab(!h2f_AWSIZE_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aligned_address_bits[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aligned_address_bits[3] .extended_lut = "off";
defparam \aligned_address_bits[3] .lut_mask = 64'h4444444444444444;
defparam \aligned_address_bits[3] .shared_arith = "off";

cyclonev_lcell_comb \aligned_address_bits[1] (
	.dataa(!h2f_AWADDR_1),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aligned_address_bits[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aligned_address_bits[1] .extended_lut = "off";
defparam \aligned_address_bits[1] .lut_mask = 64'h4040404040404040;
defparam \aligned_address_bits[1] .shared_arith = "off";

cyclonev_lcell_comb \Add0~109 (
	.dataa(!sop_enable),
	.datab(!address_burst_0),
	.datac(!h2f_AWADDR_0),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!Decoder01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(\Add0~110 ),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h0000EEE4000000FF;
defparam \Add0~109 .shared_arith = "off";

cyclonev_lcell_comb \Add0~105 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!address_burst_1),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!\aligned_address_bits[1]~combout ),
	.datag(gnd),
	.cin(\Add0~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h0000FA50000000FF;
defparam \Add0~105 .shared_arith = "off";

cyclonev_lcell_comb \Add0~89 (
	.dataa(!sop_enable),
	.datab(!address_burst_2),
	.datac(!h2f_AWADDR_2),
	.datad(!Decoder04),
	.datae(gnd),
	.dataf(!LessThan2),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h0000E4EE000000FF;
defparam \Add0~89 .shared_arith = "off";

cyclonev_lcell_comb \Add0~93 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!address_burst_3),
	.datad(!Decoder05),
	.datae(gnd),
	.dataf(!\aligned_address_bits[3]~combout ),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h0000FA50000000FF;
defparam \Add0~93 .shared_arith = "off";

cyclonev_lcell_comb \Add0~97 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_4),
	.datad(!Decoder06),
	.datae(gnd),
	.dataf(!address_burst_4),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~97 .shared_arith = "off";

cyclonev_lcell_comb \Add0~101 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_5),
	.datad(!Decoder07),
	.datae(gnd),
	.dataf(!address_burst_5),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~101 .shared_arith = "off";

cyclonev_lcell_comb \Add0~81 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_6),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!address_burst_6),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~81 .shared_arith = "off";

cyclonev_lcell_comb \Add0~73 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_7),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!address_burst_7),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~73 .shared_arith = "off";

cyclonev_lcell_comb \Add0~85 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_8),
	.datad(!address_burst_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~85 .shared_arith = "off";

cyclonev_lcell_comb \Add0~77 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_9),
	.datad(!address_burst_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~77 .shared_arith = "off";

cyclonev_lcell_comb \Add0~65 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_10),
	.datad(!address_burst_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~65 .shared_arith = "off";

cyclonev_lcell_comb \Add0~69 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_11),
	.datad(!address_burst_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~69 .shared_arith = "off";

cyclonev_lcell_comb \Add0~57 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_12),
	.datad(!address_burst_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~57 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_13),
	.datad(!address_burst_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~61 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_14),
	.datad(!address_burst_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~61 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_15),
	.datad(!address_burst_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_16),
	.datad(!address_burst_16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_17),
	.datad(!address_burst_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_18),
	.datad(!address_burst_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~45 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_19),
	.datad(!address_burst_19),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_20),
	.datad(!address_burst_20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_21),
	.datad(!address_burst_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_22),
	.datad(!address_burst_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_23),
	.datad(!address_burst_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_24),
	.datad(!address_burst_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[24]~2 (
	.dataa(!h2f_AWADDR_24),
	.datab(!sop_enable),
	.datac(!address_burst_24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[24]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[24]~2 .extended_lut = "off";
defparam \out_data[24]~2 .lut_mask = 64'h4747474747474747;
defparam \out_data[24]~2 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_25),
	.datad(!address_burst_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \out_data[25]~3 (
	.dataa(!h2f_AWADDR_25),
	.datab(!sop_enable),
	.datac(!address_burst_25),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[25]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[25]~3 .extended_lut = "off";
defparam \out_data[25]~3 .lut_mask = 64'h4747474747474747;
defparam \out_data[25]~3 .shared_arith = "off";

cyclonev_lcell_comb \out_data[23]~4 (
	.dataa(!h2f_AWADDR_23),
	.datab(!sop_enable),
	.datac(!address_burst_23),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[23]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[23]~4 .extended_lut = "off";
defparam \out_data[23]~4 .lut_mask = 64'h4747474747474747;
defparam \out_data[23]~4 .shared_arith = "off";

cyclonev_lcell_comb \out_data[13]~5 (
	.dataa(!h2f_AWADDR_13),
	.datab(!sop_enable),
	.datac(!address_burst_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[13]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[13]~5 .extended_lut = "off";
defparam \out_data[13]~5 .lut_mask = 64'h4747474747474747;
defparam \out_data[13]~5 .shared_arith = "off";

cyclonev_lcell_comb \out_data[21]~6 (
	.dataa(!h2f_AWADDR_21),
	.datab(!sop_enable),
	.datac(!address_burst_21),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[21]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[21]~6 .extended_lut = "off";
defparam \out_data[21]~6 .lut_mask = 64'h4747474747474747;
defparam \out_data[21]~6 .shared_arith = "off";

cyclonev_lcell_comb \out_data[22]~7 (
	.dataa(!h2f_AWADDR_22),
	.datab(!sop_enable),
	.datac(!address_burst_22),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[22]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[22]~7 .extended_lut = "off";
defparam \out_data[22]~7 .lut_mask = 64'h4747474747474747;
defparam \out_data[22]~7 .shared_arith = "off";

cyclonev_lcell_comb \out_data[19]~8 (
	.dataa(!h2f_AWADDR_19),
	.datab(!sop_enable),
	.datac(!address_burst_19),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[19]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[19]~8 .extended_lut = "off";
defparam \out_data[19]~8 .lut_mask = 64'h4747474747474747;
defparam \out_data[19]~8 .shared_arith = "off";

cyclonev_lcell_comb \out_data[20]~9 (
	.dataa(!h2f_AWADDR_20),
	.datab(!sop_enable),
	.datac(!address_burst_20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[20]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[20]~9 .extended_lut = "off";
defparam \out_data[20]~9 .lut_mask = 64'h4747474747474747;
defparam \out_data[20]~9 .shared_arith = "off";

cyclonev_lcell_comb \out_data[15]~10 (
	.dataa(!h2f_AWADDR_15),
	.datab(!sop_enable),
	.datac(!address_burst_15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[15]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[15]~10 .extended_lut = "off";
defparam \out_data[15]~10 .lut_mask = 64'h4747474747474747;
defparam \out_data[15]~10 .shared_arith = "off";

cyclonev_lcell_comb \out_data[16]~11 (
	.dataa(!h2f_AWADDR_16),
	.datab(!sop_enable),
	.datac(!address_burst_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[16]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[16]~11 .extended_lut = "off";
defparam \out_data[16]~11 .lut_mask = 64'h4747474747474747;
defparam \out_data[16]~11 .shared_arith = "off";

cyclonev_lcell_comb \out_data[17]~12 (
	.dataa(!h2f_AWADDR_17),
	.datab(!sop_enable),
	.datac(!address_burst_17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[17]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[17]~12 .extended_lut = "off";
defparam \out_data[17]~12 .lut_mask = 64'h4747474747474747;
defparam \out_data[17]~12 .shared_arith = "off";

cyclonev_lcell_comb \out_data[18]~13 (
	.dataa(!h2f_AWADDR_18),
	.datab(!sop_enable),
	.datac(!address_burst_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[18]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[18]~13 .extended_lut = "off";
defparam \out_data[18]~13 .lut_mask = 64'h4747474747474747;
defparam \out_data[18]~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~49 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_26),
	.datad(!address_burst_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~49 .shared_arith = "off";

cyclonev_lcell_comb \out_data[26]~14 (
	.dataa(!h2f_AWADDR_26),
	.datab(!sop_enable),
	.datac(!address_burst_26),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[26]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[26]~14 .extended_lut = "off";
defparam \out_data[26]~14 .lut_mask = 64'h4747474747474747;
defparam \out_data[26]~14 .shared_arith = "off";

cyclonev_lcell_comb \Add0~53 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_27),
	.datad(!address_burst_27),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~53 .shared_arith = "off";

cyclonev_lcell_comb \out_data[27]~15 (
	.dataa(!h2f_AWADDR_27),
	.datab(!sop_enable),
	.datac(!address_burst_27),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[27]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[27]~15 .extended_lut = "off";
defparam \out_data[27]~15 .lut_mask = 64'h4747474747474747;
defparam \out_data[27]~15 .shared_arith = "off";

cyclonev_lcell_comb \out_data[12]~16 (
	.dataa(!h2f_AWADDR_12),
	.datab(!sop_enable),
	.datac(!address_burst_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[12]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[12]~16 .extended_lut = "off";
defparam \out_data[12]~16 .lut_mask = 64'h4747474747474747;
defparam \out_data[12]~16 .shared_arith = "off";

cyclonev_lcell_comb \out_data[14]~17 (
	.dataa(!h2f_AWADDR_14),
	.datab(!sop_enable),
	.datac(!address_burst_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[14]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[14]~17 .extended_lut = "off";
defparam \out_data[14]~17 .lut_mask = 64'h4747474747474747;
defparam \out_data[14]~17 .shared_arith = "off";

cyclonev_lcell_comb \out_data[10]~18 (
	.dataa(!h2f_AWADDR_10),
	.datab(!sop_enable),
	.datac(!address_burst_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[10]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[10]~18 .extended_lut = "off";
defparam \out_data[10]~18 .lut_mask = 64'h4747474747474747;
defparam \out_data[10]~18 .shared_arith = "off";

cyclonev_lcell_comb \out_data[11]~19 (
	.dataa(!h2f_AWADDR_11),
	.datab(!sop_enable),
	.datac(!address_burst_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[11]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[11]~19 .extended_lut = "off";
defparam \out_data[11]~19 .lut_mask = 64'h4747474747474747;
defparam \out_data[11]~19 .shared_arith = "off";

cyclonev_lcell_comb \Add1~29 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!address_burst_0),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!h2f_AWADDR_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~29_sumout ),
	.cout(\Add1~30 ),
	.shareout());
defparam \Add1~29 .extended_lut = "off";
defparam \Add1~29 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~29 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!address_burst_1),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!h2f_AWADDR_1),
	.datag(gnd),
	.cin(\Add1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~25 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!address_burst_2),
	.datad(!Decoder04),
	.datae(gnd),
	.dataf(!h2f_AWADDR_2),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!address_burst_3),
	.datad(!Decoder05),
	.datae(gnd),
	.dataf(!h2f_AWADDR_3),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_4),
	.datad(!Decoder06),
	.datae(gnd),
	.dataf(!address_burst_4),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_5),
	.datad(!Decoder07),
	.datae(gnd),
	.dataf(!address_burst_5),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_6),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!address_burst_6),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_AWADDR_7),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!address_burst_7),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector22~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!out_data_7),
	.datad(!Add11),
	.datae(!\Add1~1_sumout ),
	.dataf(!\Add0~73_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector22~0 .extended_lut = "off";
defparam \Selector22~0 .lut_mask = 64'h0A080A2A5F5D5F7F;
defparam \Selector22~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector23~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!out_data_6),
	.datad(!LessThan16),
	.datae(!\Add1~5_sumout ),
	.dataf(!\Add0~81_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector23~0 .extended_lut = "off";
defparam \Selector23~0 .lut_mask = 64'h080A2A0A5D5F7F5F;
defparam \Selector23~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector27~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!out_data_2),
	.datad(!LessThan12),
	.datae(!\Add1~9_sumout ),
	.dataf(!\Add0~89_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~0 .extended_lut = "off";
defparam \Selector27~0 .lut_mask = 64'h080A2A0A5D5F7F5F;
defparam \Selector27~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~1 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!out_data_3),
	.datad(!Selector26),
	.datae(!\Add1~13_sumout ),
	.dataf(!\Add0~93_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~1 .extended_lut = "off";
defparam \Selector26~1 .lut_mask = 64'h080A2A0A5D5F7F5F;
defparam \Selector26~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector25~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!out_data_4),
	.datad(!\Add1~17_sumout ),
	.datae(!LessThan14),
	.dataf(!\Add0~97_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~0 .extended_lut = "off";
defparam \Selector25~0 .lut_mask = 64'h082A0A0A5D7F5F5F;
defparam \Selector25~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector24~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!out_data_5),
	.datad(!LessThan15),
	.datae(!\Add1~21_sumout ),
	.dataf(!\Add0~101_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~0 .extended_lut = "off";
defparam \Selector24~0 .lut_mask = 64'h080A2A0A5D5F7F5F;
defparam \Selector24~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!LessThan11),
	.datad(!out_data_1),
	.datae(!\Add1~25_sumout ),
	.dataf(!\Add0~105_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~0 .extended_lut = "off";
defparam \Selector28~0 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector28~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector29~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!LessThan10),
	.datad(!out_data_0),
	.datae(!\Add1~29_sumout ),
	.dataf(!\Add0~109_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector29~0 .extended_lut = "off";
defparam \Selector29~0 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector29~0 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_burst_adapter (
	h2f_AWBURST_0,
	h2f_AWBURST_1,
	outclk_wire_0,
	Add4,
	Add41,
	out_data_37,
	Mux4,
	Mux5,
	Mux6,
	Mux7,
	Mux8,
	Mux9,
	Mux10,
	Mux11,
	Mux12,
	Mux13,
	Mux14,
	Mux15,
	Mux16,
	Mux17,
	Mux18,
	Mux19,
	Mux20,
	Mux21,
	Mux22,
	Mux23,
	Mux24,
	Mux25,
	Mux26,
	Mux27,
	Mux28,
	Mux29,
	Mux30,
	Mux31,
	Mux32,
	Mux33,
	Mux34,
	Mux35,
	Mux3,
	Mux2,
	Mux1,
	Mux0,
	in_ready_hold,
	Equal0,
	Equal01,
	Equal02,
	nxt_in_ready,
	out_valid_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wrfull,
	wrfull1,
	wrfull2,
	mem_used_1,
	load_next_out_cmd,
	saved_grant_0,
	in_data_reg_68,
	nxt_uncomp_subburst_byte_cnt,
	in_data_reg_0,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	r_sync_rst,
	LessThan12,
	Selector26,
	src0_valid,
	in_eop_reg,
	wrfull3,
	int_output_sel_0,
	int_output_sel_1,
	cp_ready,
	src_payload,
	src_payload1,
	src_payload2,
	in_data_reg_122,
	in_data_reg_123,
	in_data_reg_124,
	in_data_reg_90,
	in_data_reg_91,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	in_data_reg_104,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	Selector7,
	Selector8,
	out_endofpacket,
	nxt_in_ready1,
	nxt_in_ready2,
	out_data_90,
	out_data_91,
	out_burstwrap_reg_2,
	out_burstwrap_reg_3,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	out_addr_reg_1,
	out_data_36,
	out_burstwrap_reg_1,
	out_addr_reg_0,
	src_payload15,
	out_burstwrap_reg_0)/* synthesis synthesis_greybox=0 */;
input 	h2f_AWBURST_0;
input 	h2f_AWBURST_1;
input 	outclk_wire_0;
input 	Add4;
input 	Add41;
input 	out_data_37;
input 	Mux4;
input 	Mux5;
input 	Mux6;
input 	Mux7;
input 	Mux8;
input 	Mux9;
input 	Mux10;
input 	Mux11;
input 	Mux12;
input 	Mux13;
input 	Mux14;
input 	Mux15;
input 	Mux16;
input 	Mux17;
input 	Mux18;
input 	Mux19;
input 	Mux20;
input 	Mux21;
input 	Mux22;
input 	Mux23;
input 	Mux24;
input 	Mux25;
input 	Mux26;
input 	Mux27;
input 	Mux28;
input 	Mux29;
input 	Mux30;
input 	Mux31;
input 	Mux32;
input 	Mux33;
input 	Mux34;
input 	Mux35;
input 	Mux3;
input 	Mux2;
input 	Mux1;
input 	Mux0;
input 	in_ready_hold;
input 	Equal0;
input 	Equal01;
input 	Equal02;
output 	nxt_in_ready;
output 	out_valid_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
input 	WideOr0;
input 	wrfull;
input 	wrfull1;
input 	wrfull2;
input 	mem_used_1;
output 	load_next_out_cmd;
input 	saved_grant_0;
output 	in_data_reg_68;
output 	nxt_uncomp_subburst_byte_cnt;
output 	in_data_reg_0;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
input 	r_sync_rst;
input 	LessThan12;
input 	Selector26;
input 	src0_valid;
output 	in_eop_reg;
input 	wrfull3;
input 	int_output_sel_0;
input 	int_output_sel_1;
input 	cp_ready;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
output 	in_data_reg_122;
output 	in_data_reg_123;
output 	in_data_reg_124;
output 	in_data_reg_90;
output 	in_data_reg_91;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_3;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
output 	in_data_reg_104;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
input 	Selector7;
input 	Selector8;
input 	out_endofpacket;
output 	nxt_in_ready1;
output 	nxt_in_ready2;
input 	out_data_90;
input 	out_data_91;
output 	out_burstwrap_reg_2;
output 	out_burstwrap_reg_3;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
output 	out_addr_reg_1;
input 	out_data_36;
output 	out_burstwrap_reg_1;
output 	out_addr_reg_0;
input 	src_payload15;
output 	out_burstwrap_reg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altera_merlin_burst_adapter_13_1 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_AWBURST_0(h2f_AWBURST_0),
	.h2f_AWBURST_1(h2f_AWBURST_1),
	.outclk_wire_0(outclk_wire_0),
	.Add4(Add4),
	.Add41(Add41),
	.out_data_37(out_data_37),
	.sink0_data({src_payload2,src_payload,src_payload1,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload14,src_payload13,src_payload12,src_payload11,src_payload10,src_payload9,src_payload8,src_payload7,src_payload6,src_payload5,src_payload4,src_payload3,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,out_data_91,
out_data_90,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload15,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux0,Mux1,Mux2,Mux3,Mux4,Mux5,Mux6,Mux7,Mux8,Mux9,Mux10,Mux11,Mux12,Mux13,
Mux14,Mux15,Mux16,Mux17,Mux18,Mux19,Mux20,Mux21,Mux22,Mux23,Mux24,Mux25,Mux26,Mux27,Mux28,Mux29,Mux30,Mux31,Mux32,Mux33,Mux34,Mux35}),
	.in_ready_hold(in_ready_hold),
	.Equal0(Equal0),
	.Equal01(Equal01),
	.Equal02(Equal02),
	.nxt_in_ready(nxt_in_ready),
	.out_valid_reg1(out_valid_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.WideOr0(WideOr0),
	.wrfull(wrfull),
	.wrfull1(wrfull1),
	.wrfull2(wrfull2),
	.mem_used_1(mem_used_1),
	.load_next_out_cmd1(load_next_out_cmd),
	.in_data_reg_68(in_data_reg_68),
	.nxt_uncomp_subburst_byte_cnt(nxt_uncomp_subburst_byte_cnt),
	.in_data_reg_0(in_data_reg_0),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_24(in_data_reg_24),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_31(in_data_reg_31),
	.r_sync_rst(r_sync_rst),
	.LessThan12(LessThan12),
	.Selector26(Selector26),
	.src0_valid(src0_valid),
	.in_eop_reg1(in_eop_reg),
	.wrfull3(wrfull3),
	.int_output_sel_0(int_output_sel_0),
	.int_output_sel_1(int_output_sel_1),
	.cp_ready(cp_ready),
	.in_data_reg_122(in_data_reg_122),
	.in_data_reg_123(in_data_reg_123),
	.in_data_reg_124(in_data_reg_124),
	.in_data_reg_90(in_data_reg_90),
	.in_data_reg_91(in_data_reg_91),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.in_data_reg_101(in_data_reg_101),
	.in_data_reg_102(in_data_reg_102),
	.in_data_reg_103(in_data_reg_103),
	.in_data_reg_104(in_data_reg_104),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.Selector7(Selector7),
	.Selector8(Selector8),
	.sink0_endofpacket(out_endofpacket),
	.nxt_in_ready1(nxt_in_ready1),
	.nxt_in_ready2(nxt_in_ready2),
	.out_burstwrap_reg_2(out_burstwrap_reg_2),
	.out_burstwrap_reg_3(out_burstwrap_reg_3),
	.out_addr_reg_1(out_addr_reg_1),
	.out_data_36(out_data_36),
	.out_burstwrap_reg_1(out_burstwrap_reg_1),
	.out_addr_reg_0(out_addr_reg_0),
	.out_burstwrap_reg_0(out_burstwrap_reg_0));

endmodule

module Computer_System_altera_merlin_burst_adapter_13_1 (
	h2f_AWBURST_0,
	h2f_AWBURST_1,
	outclk_wire_0,
	Add4,
	Add41,
	out_data_37,
	sink0_data,
	in_ready_hold,
	Equal0,
	Equal01,
	Equal02,
	nxt_in_ready,
	out_valid_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wrfull,
	wrfull1,
	wrfull2,
	mem_used_1,
	load_next_out_cmd1,
	in_data_reg_68,
	nxt_uncomp_subburst_byte_cnt,
	in_data_reg_0,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	r_sync_rst,
	LessThan12,
	Selector26,
	src0_valid,
	in_eop_reg1,
	wrfull3,
	int_output_sel_0,
	int_output_sel_1,
	cp_ready,
	in_data_reg_122,
	in_data_reg_123,
	in_data_reg_124,
	in_data_reg_90,
	in_data_reg_91,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	in_data_reg_104,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	Selector7,
	Selector8,
	sink0_endofpacket,
	nxt_in_ready1,
	nxt_in_ready2,
	out_burstwrap_reg_2,
	out_burstwrap_reg_3,
	out_addr_reg_1,
	out_data_36,
	out_burstwrap_reg_1,
	out_addr_reg_0,
	out_burstwrap_reg_0)/* synthesis synthesis_greybox=0 */;
input 	h2f_AWBURST_0;
input 	h2f_AWBURST_1;
input 	outclk_wire_0;
input 	Add4;
input 	Add41;
input 	out_data_37;
input 	[124:0] sink0_data;
input 	in_ready_hold;
input 	Equal0;
input 	Equal01;
input 	Equal02;
output 	nxt_in_ready;
output 	out_valid_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
input 	WideOr0;
input 	wrfull;
input 	wrfull1;
input 	wrfull2;
input 	mem_used_1;
output 	load_next_out_cmd1;
output 	in_data_reg_68;
output 	nxt_uncomp_subburst_byte_cnt;
output 	in_data_reg_0;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
input 	r_sync_rst;
input 	LessThan12;
input 	Selector26;
input 	src0_valid;
output 	in_eop_reg1;
input 	wrfull3;
input 	int_output_sel_0;
input 	int_output_sel_1;
input 	cp_ready;
output 	in_data_reg_122;
output 	in_data_reg_123;
output 	in_data_reg_124;
output 	in_data_reg_90;
output 	in_data_reg_91;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_3;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
output 	in_data_reg_104;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
input 	Selector7;
input 	Selector8;
input 	sink0_endofpacket;
output 	nxt_in_ready1;
output 	nxt_in_ready2;
output 	out_burstwrap_reg_2;
output 	out_burstwrap_reg_3;
output 	out_addr_reg_1;
input 	out_data_36;
output 	out_burstwrap_reg_1;
output 	out_addr_reg_0;
output 	out_burstwrap_reg_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \in_valid~0_combout ;
wire \Selector0~0_combout ;
wire \state.ST_IDLE~q ;
wire \new_burst_reg~q ;
wire \nxt_uncomp_subburst_byte_cnt[2]~6_combout ;
wire \out_uncomp_byte_cnt_reg[2]~q ;
wire \Add4~1_sumout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~7_combout ;
wire \out_uncomp_byte_cnt_reg[3]~q ;
wire \Add4~2 ;
wire \Add4~3 ;
wire \Add4~5_sumout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~3_combout ;
wire \out_uncomp_byte_cnt_reg[4]~q ;
wire \Add4~6 ;
wire \Add4~7 ;
wire \Add4~9_sumout ;
wire \Add4~10 ;
wire \Add4~11 ;
wire \Add4~13_sumout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~1_combout ;
wire \out_uncomp_byte_cnt_reg[5]~q ;
wire \Add4~14 ;
wire \Add4~15 ;
wire \Add4~17_sumout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~2_combout ;
wire \out_uncomp_byte_cnt_reg[6]~q ;
wire \WideOr0~4_combout ;
wire \WideOr0~0_combout ;
wire \Add4~18 ;
wire \Add4~19 ;
wire \Add4~25_sumout ;
wire \nxt_uncomp_subburst_byte_cnt[7]~5_combout ;
wire \out_uncomp_byte_cnt_reg[7]~q ;
wire \Add4~26 ;
wire \Add4~27 ;
wire \Add4~21_sumout ;
wire \nxt_uncomp_subburst_byte_cnt[8]~4_combout ;
wire \out_uncomp_byte_cnt_reg[8]~q ;
wire \WideOr0~5_combout ;
wire \WideOr0~1_combout ;
wire \WideOr0~2_combout ;
wire \WideOr0~3_combout ;
wire \Selector2~0_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector3~1_combout ;
wire \Selector3~2_combout ;
wire \Selector3~0_combout ;
wire \state.ST_UNCOMP_WR_SUBBURST~q ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \nxt_out_burstwrap[2]~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_out_burstwrap[2]~1_combout ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \nxt_out_burstwrap[0]~5_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_out_burstwrap[0]~6_combout ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_out_burstwrap[1]~4_combout ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \out_addr_reg~0_combout ;
wire \d0_int_nxt_addr[1]~2_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[2]~0_combout ;
wire \nxt_out_burstwrap[3]~2_combout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_out_burstwrap[3]~3_combout ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[3]~1_combout ;
wire \out_addr_reg~1_combout ;
wire \out_addr_reg~2_combout ;


Computer_System_altera_merlin_address_alignment_1 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.in_data_reg_90(in_data_reg_90),
	.in_data_reg_91(in_data_reg_91),
	.out_data_90(sink0_data[90]),
	.out_data_91(sink0_data[91]),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\state.ST_UNCOMP_WR_SUBBURST~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h8888888888888888;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(outclk_wire_0),
	.d(\in_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!WideOr0),
	.datac(!wrfull),
	.datad(!wrfull1),
	.datae(!wrfull2),
	.dataf(!mem_used_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(load_next_out_cmd1),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBFFFBAAAAAAAA;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \in_data_reg[68] (
	.clk(outclk_wire_0),
	.d(sink0_data[68]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_68),
	.prn(vcc));
defparam \in_data_reg[68] .is_wysiwyg = "true";
defparam \in_data_reg[68] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_uncomp_subburst_byte_cnt),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h4444444444444444;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \in_data_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_1),
	.prn(vcc));
defparam \in_data_reg[1] .is_wysiwyg = "true";
defparam \in_data_reg[1] .power_up = "low";

dffeas \in_data_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_2),
	.prn(vcc));
defparam \in_data_reg[2] .is_wysiwyg = "true";
defparam \in_data_reg[2] .power_up = "low";

dffeas \in_data_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_3),
	.prn(vcc));
defparam \in_data_reg[3] .is_wysiwyg = "true";
defparam \in_data_reg[3] .power_up = "low";

dffeas \in_data_reg[4] (
	.clk(outclk_wire_0),
	.d(sink0_data[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_4),
	.prn(vcc));
defparam \in_data_reg[4] .is_wysiwyg = "true";
defparam \in_data_reg[4] .power_up = "low";

dffeas \in_data_reg[5] (
	.clk(outclk_wire_0),
	.d(sink0_data[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_5),
	.prn(vcc));
defparam \in_data_reg[5] .is_wysiwyg = "true";
defparam \in_data_reg[5] .power_up = "low";

dffeas \in_data_reg[6] (
	.clk(outclk_wire_0),
	.d(sink0_data[6]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_6),
	.prn(vcc));
defparam \in_data_reg[6] .is_wysiwyg = "true";
defparam \in_data_reg[6] .power_up = "low";

dffeas \in_data_reg[7] (
	.clk(outclk_wire_0),
	.d(sink0_data[7]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_7),
	.prn(vcc));
defparam \in_data_reg[7] .is_wysiwyg = "true";
defparam \in_data_reg[7] .power_up = "low";

dffeas \in_data_reg[8] (
	.clk(outclk_wire_0),
	.d(sink0_data[8]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_8),
	.prn(vcc));
defparam \in_data_reg[8] .is_wysiwyg = "true";
defparam \in_data_reg[8] .power_up = "low";

dffeas \in_data_reg[9] (
	.clk(outclk_wire_0),
	.d(sink0_data[9]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_9),
	.prn(vcc));
defparam \in_data_reg[9] .is_wysiwyg = "true";
defparam \in_data_reg[9] .power_up = "low";

dffeas \in_data_reg[10] (
	.clk(outclk_wire_0),
	.d(sink0_data[10]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_10),
	.prn(vcc));
defparam \in_data_reg[10] .is_wysiwyg = "true";
defparam \in_data_reg[10] .power_up = "low";

dffeas \in_data_reg[11] (
	.clk(outclk_wire_0),
	.d(sink0_data[11]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_11),
	.prn(vcc));
defparam \in_data_reg[11] .is_wysiwyg = "true";
defparam \in_data_reg[11] .power_up = "low";

dffeas \in_data_reg[12] (
	.clk(outclk_wire_0),
	.d(sink0_data[12]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_12),
	.prn(vcc));
defparam \in_data_reg[12] .is_wysiwyg = "true";
defparam \in_data_reg[12] .power_up = "low";

dffeas \in_data_reg[13] (
	.clk(outclk_wire_0),
	.d(sink0_data[13]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_13),
	.prn(vcc));
defparam \in_data_reg[13] .is_wysiwyg = "true";
defparam \in_data_reg[13] .power_up = "low";

dffeas \in_data_reg[14] (
	.clk(outclk_wire_0),
	.d(sink0_data[14]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_14),
	.prn(vcc));
defparam \in_data_reg[14] .is_wysiwyg = "true";
defparam \in_data_reg[14] .power_up = "low";

dffeas \in_data_reg[15] (
	.clk(outclk_wire_0),
	.d(sink0_data[15]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_15),
	.prn(vcc));
defparam \in_data_reg[15] .is_wysiwyg = "true";
defparam \in_data_reg[15] .power_up = "low";

dffeas \in_data_reg[16] (
	.clk(outclk_wire_0),
	.d(sink0_data[16]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_16),
	.prn(vcc));
defparam \in_data_reg[16] .is_wysiwyg = "true";
defparam \in_data_reg[16] .power_up = "low";

dffeas \in_data_reg[17] (
	.clk(outclk_wire_0),
	.d(sink0_data[17]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_17),
	.prn(vcc));
defparam \in_data_reg[17] .is_wysiwyg = "true";
defparam \in_data_reg[17] .power_up = "low";

dffeas \in_data_reg[18] (
	.clk(outclk_wire_0),
	.d(sink0_data[18]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_18),
	.prn(vcc));
defparam \in_data_reg[18] .is_wysiwyg = "true";
defparam \in_data_reg[18] .power_up = "low";

dffeas \in_data_reg[19] (
	.clk(outclk_wire_0),
	.d(sink0_data[19]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_19),
	.prn(vcc));
defparam \in_data_reg[19] .is_wysiwyg = "true";
defparam \in_data_reg[19] .power_up = "low";

dffeas \in_data_reg[20] (
	.clk(outclk_wire_0),
	.d(sink0_data[20]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_20),
	.prn(vcc));
defparam \in_data_reg[20] .is_wysiwyg = "true";
defparam \in_data_reg[20] .power_up = "low";

dffeas \in_data_reg[21] (
	.clk(outclk_wire_0),
	.d(sink0_data[21]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_21),
	.prn(vcc));
defparam \in_data_reg[21] .is_wysiwyg = "true";
defparam \in_data_reg[21] .power_up = "low";

dffeas \in_data_reg[22] (
	.clk(outclk_wire_0),
	.d(sink0_data[22]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_22),
	.prn(vcc));
defparam \in_data_reg[22] .is_wysiwyg = "true";
defparam \in_data_reg[22] .power_up = "low";

dffeas \in_data_reg[23] (
	.clk(outclk_wire_0),
	.d(sink0_data[23]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_23),
	.prn(vcc));
defparam \in_data_reg[23] .is_wysiwyg = "true";
defparam \in_data_reg[23] .power_up = "low";

dffeas \in_data_reg[24] (
	.clk(outclk_wire_0),
	.d(sink0_data[24]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_24),
	.prn(vcc));
defparam \in_data_reg[24] .is_wysiwyg = "true";
defparam \in_data_reg[24] .power_up = "low";

dffeas \in_data_reg[25] (
	.clk(outclk_wire_0),
	.d(sink0_data[25]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_25),
	.prn(vcc));
defparam \in_data_reg[25] .is_wysiwyg = "true";
defparam \in_data_reg[25] .power_up = "low";

dffeas \in_data_reg[26] (
	.clk(outclk_wire_0),
	.d(sink0_data[26]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_26),
	.prn(vcc));
defparam \in_data_reg[26] .is_wysiwyg = "true";
defparam \in_data_reg[26] .power_up = "low";

dffeas \in_data_reg[27] (
	.clk(outclk_wire_0),
	.d(sink0_data[27]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_27),
	.prn(vcc));
defparam \in_data_reg[27] .is_wysiwyg = "true";
defparam \in_data_reg[27] .power_up = "low";

dffeas \in_data_reg[28] (
	.clk(outclk_wire_0),
	.d(sink0_data[28]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_28),
	.prn(vcc));
defparam \in_data_reg[28] .is_wysiwyg = "true";
defparam \in_data_reg[28] .power_up = "low";

dffeas \in_data_reg[29] (
	.clk(outclk_wire_0),
	.d(sink0_data[29]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_29),
	.prn(vcc));
defparam \in_data_reg[29] .is_wysiwyg = "true";
defparam \in_data_reg[29] .power_up = "low";

dffeas \in_data_reg[30] (
	.clk(outclk_wire_0),
	.d(sink0_data[30]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_30),
	.prn(vcc));
defparam \in_data_reg[30] .is_wysiwyg = "true";
defparam \in_data_reg[30] .power_up = "low";

dffeas \in_data_reg[31] (
	.clk(outclk_wire_0),
	.d(sink0_data[31]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_31),
	.prn(vcc));
defparam \in_data_reg[31] .is_wysiwyg = "true";
defparam \in_data_reg[31] .power_up = "low";

dffeas in_eop_reg(
	.clk(outclk_wire_0),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_eop_reg1),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

dffeas \in_data_reg[122] (
	.clk(outclk_wire_0),
	.d(sink0_data[122]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_122),
	.prn(vcc));
defparam \in_data_reg[122] .is_wysiwyg = "true";
defparam \in_data_reg[122] .power_up = "low";

dffeas \in_data_reg[123] (
	.clk(outclk_wire_0),
	.d(sink0_data[123]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_123),
	.prn(vcc));
defparam \in_data_reg[123] .is_wysiwyg = "true";
defparam \in_data_reg[123] .power_up = "low";

dffeas \in_data_reg[124] (
	.clk(outclk_wire_0),
	.d(sink0_data[124]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_124),
	.prn(vcc));
defparam \in_data_reg[124] .is_wysiwyg = "true";
defparam \in_data_reg[124] .power_up = "low";

dffeas \in_data_reg[90] (
	.clk(outclk_wire_0),
	.d(sink0_data[90]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_90),
	.prn(vcc));
defparam \in_data_reg[90] .is_wysiwyg = "true";
defparam \in_data_reg[90] .power_up = "low";

dffeas \in_data_reg[91] (
	.clk(outclk_wire_0),
	.d(sink0_data[91]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_91),
	.prn(vcc));
defparam \in_data_reg[91] .is_wysiwyg = "true";
defparam \in_data_reg[91] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[2]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[3]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \in_data_reg[101] (
	.clk(outclk_wire_0),
	.d(sink0_data[101]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_101),
	.prn(vcc));
defparam \in_data_reg[101] .is_wysiwyg = "true";
defparam \in_data_reg[101] .power_up = "low";

dffeas \in_data_reg[102] (
	.clk(outclk_wire_0),
	.d(sink0_data[102]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_102),
	.prn(vcc));
defparam \in_data_reg[102] .is_wysiwyg = "true";
defparam \in_data_reg[102] .power_up = "low";

dffeas \in_data_reg[103] (
	.clk(outclk_wire_0),
	.d(sink0_data[103]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_103),
	.prn(vcc));
defparam \in_data_reg[103] .is_wysiwyg = "true";
defparam \in_data_reg[103] .power_up = "low";

dffeas \in_data_reg[104] (
	.clk(outclk_wire_0),
	.d(sink0_data[104]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_104),
	.prn(vcc));
defparam \in_data_reg[104] .is_wysiwyg = "true";
defparam \in_data_reg[104] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(outclk_wire_0),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(outclk_wire_0),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(outclk_wire_0),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(outclk_wire_0),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(outclk_wire_0),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(outclk_wire_0),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(outclk_wire_0),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(outclk_wire_0),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!in_ready_hold),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!\state.ST_UNCOMP_WR_SUBBURST~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h4040404040404040;
defparam \nxt_in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~2 (
	.dataa(!nxt_in_ready),
	.datab(!out_valid_reg1),
	.datac(!WideOr0),
	.datad(!wrfull3),
	.datae(!wrfull2),
	.dataf(!mem_used_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~2 .extended_lut = "off";
defparam \nxt_in_ready~2 .lut_mask = 64'h8A8AAA8A88888888;
defparam \nxt_in_ready~2 .shared_arith = "off";

dffeas \out_burstwrap_reg[2] (
	.clk(outclk_wire_0),
	.d(\nxt_out_burstwrap[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(out_burstwrap_reg_2),
	.prn(vcc));
defparam \out_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \out_burstwrap_reg[2] .power_up = "low";

dffeas \out_burstwrap_reg[3] (
	.clk(outclk_wire_0),
	.d(\nxt_out_burstwrap[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(out_burstwrap_reg_3),
	.prn(vcc));
defparam \out_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \out_burstwrap_reg[3] .power_up = "low";

dffeas \out_addr_reg[1] (
	.clk(outclk_wire_0),
	.d(\out_addr_reg~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(out_addr_reg_1),
	.prn(vcc));
defparam \out_addr_reg[1] .is_wysiwyg = "true";
defparam \out_addr_reg[1] .power_up = "low";

dffeas \out_burstwrap_reg[1] (
	.clk(outclk_wire_0),
	.d(\nxt_out_burstwrap[1]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(out_burstwrap_reg_1),
	.prn(vcc));
defparam \out_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \out_burstwrap_reg[1] .power_up = "low";

dffeas \out_addr_reg[0] (
	.clk(outclk_wire_0),
	.d(\out_addr_reg~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(out_addr_reg_0),
	.prn(vcc));
defparam \out_addr_reg[0] .is_wysiwyg = "true";
defparam \out_addr_reg[0] .power_up = "low";

dffeas \out_burstwrap_reg[0] (
	.clk(outclk_wire_0),
	.d(\nxt_out_burstwrap[0]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(out_burstwrap_reg_0),
	.prn(vcc));
defparam \out_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \out_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \in_valid~0 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[68]),
	.datac(!Equal0),
	.datad(!Equal01),
	.datae(!Equal02),
	.dataf(!src0_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_valid~0 .extended_lut = "off";
defparam \in_valid~0 .lut_mask = 64'h0000000000000001;
defparam \in_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!\state.ST_IDLE~q ),
	.datab(!\in_valid~0_combout ),
	.datac(!in_eop_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h7373737373737373;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(outclk_wire_0),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

dffeas new_burst_reg(
	.clk(outclk_wire_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~6 (
	.dataa(!WideOr0),
	.datab(!wrfull3),
	.datac(!wrfull2),
	.datad(!nxt_uncomp_subburst_byte_cnt),
	.datae(!\out_uncomp_byte_cnt_reg[2]~q ),
	.dataf(!\new_burst_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~6 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~6 .lut_mask = 64'h005DFFFF0000FFA2;
defparam \nxt_uncomp_subburst_byte_cnt[2]~6 .shared_arith = "off";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(outclk_wire_0),
	.d(\Add4~1_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[2]~6_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(load_next_out_cmd1),
	.q(\out_uncomp_byte_cnt_reg[2]~q ),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

cyclonev_lcell_comb \Add4~1 (
	.dataa(!cp_ready),
	.datab(!out_valid_reg1),
	.datac(!\out_uncomp_byte_cnt_reg[2]~q ),
	.datad(!mem_used_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~1_sumout ),
	.cout(\Add4~2 ),
	.shareout(\Add4~3 ));
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h0000EFFF00001E0F;
defparam \Add4~1 .shared_arith = "on";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~7 (
	.dataa(!WideOr0),
	.datab(!wrfull3),
	.datac(!wrfull2),
	.datad(!nxt_uncomp_subburst_byte_cnt),
	.datae(!\out_uncomp_byte_cnt_reg[3]~q ),
	.dataf(!\new_burst_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~7 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~7 .lut_mask = 64'h005DFFFF0000FFA2;
defparam \nxt_uncomp_subburst_byte_cnt[3]~7 .shared_arith = "off";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(outclk_wire_0),
	.d(\Add4~5_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[3]~7_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(load_next_out_cmd1),
	.q(\out_uncomp_byte_cnt_reg[3]~q ),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\out_uncomp_byte_cnt_reg[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~2 ),
	.sharein(\Add4~3 ),
	.combout(),
	.sumout(\Add4~5_sumout ),
	.cout(\Add4~6 ),
	.shareout(\Add4~7 ));
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h00000F0F0000F0F0;
defparam \Add4~5 .shared_arith = "on";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~3 (
	.dataa(!WideOr0),
	.datab(!wrfull3),
	.datac(!wrfull2),
	.datad(!nxt_uncomp_subburst_byte_cnt),
	.datae(!\out_uncomp_byte_cnt_reg[4]~q ),
	.dataf(!\new_burst_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .lut_mask = 64'h005DFFFF0000FFA2;
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .shared_arith = "off";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(outclk_wire_0),
	.d(\Add4~9_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(load_next_out_cmd1),
	.q(\out_uncomp_byte_cnt_reg[4]~q ),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\out_uncomp_byte_cnt_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(\Add4~7 ),
	.combout(),
	.sumout(\Add4~9_sumout ),
	.cout(\Add4~10 ),
	.shareout(\Add4~11 ));
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add4~9 .shared_arith = "on";

cyclonev_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\out_uncomp_byte_cnt_reg[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(\Add4~11 ),
	.combout(),
	.sumout(\Add4~13_sumout ),
	.cout(\Add4~14 ),
	.shareout(\Add4~15 ));
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add4~13 .shared_arith = "on";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~1 (
	.dataa(!WideOr0),
	.datab(!wrfull3),
	.datac(!wrfull2),
	.datad(!nxt_uncomp_subburst_byte_cnt),
	.datae(!\out_uncomp_byte_cnt_reg[5]~q ),
	.dataf(!\new_burst_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .lut_mask = 64'h005DFFFF0000FFA2;
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .shared_arith = "off";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(outclk_wire_0),
	.d(\Add4~13_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(load_next_out_cmd1),
	.q(\out_uncomp_byte_cnt_reg[5]~q ),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\out_uncomp_byte_cnt_reg[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(\Add4~15 ),
	.combout(),
	.sumout(\Add4~17_sumout ),
	.cout(\Add4~18 ),
	.shareout(\Add4~19 ));
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add4~17 .shared_arith = "on";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~2 (
	.dataa(!WideOr0),
	.datab(!wrfull3),
	.datac(!wrfull2),
	.datad(!nxt_uncomp_subburst_byte_cnt),
	.datae(!\out_uncomp_byte_cnt_reg[6]~q ),
	.dataf(!\new_burst_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .lut_mask = 64'h005DFFFF0000FFA2;
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .shared_arith = "off";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(outclk_wire_0),
	.d(\Add4~17_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(load_next_out_cmd1),
	.q(\out_uncomp_byte_cnt_reg[6]~q ),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

cyclonev_lcell_comb \WideOr0~4 (
	.dataa(!\out_uncomp_byte_cnt_reg[5]~q ),
	.datab(!\out_uncomp_byte_cnt_reg[6]~q ),
	.datac(!\out_uncomp_byte_cnt_reg[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~4 .extended_lut = "off";
defparam \WideOr0~4 .lut_mask = 64'h8080808080808080;
defparam \WideOr0~4 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!WideOr0),
	.datab(!wrfull3),
	.datac(!wrfull2),
	.datad(!nxt_uncomp_subburst_byte_cnt),
	.datae(!\new_burst_reg~q ),
	.dataf(!\WideOr0~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hFFFFFFA2005D0000;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\out_uncomp_byte_cnt_reg[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~18 ),
	.sharein(\Add4~19 ),
	.combout(),
	.sumout(\Add4~25_sumout ),
	.cout(\Add4~26 ),
	.shareout(\Add4~27 ));
defparam \Add4~25 .extended_lut = "off";
defparam \Add4~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add4~25 .shared_arith = "on";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[7]~5 (
	.dataa(!WideOr0),
	.datab(!wrfull3),
	.datac(!wrfull2),
	.datad(!nxt_uncomp_subburst_byte_cnt),
	.datae(!\out_uncomp_byte_cnt_reg[7]~q ),
	.dataf(!\new_burst_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[7]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[7]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[7]~5 .lut_mask = 64'h005DFFFF0000FFA2;
defparam \nxt_uncomp_subburst_byte_cnt[7]~5 .shared_arith = "off";

dffeas \out_uncomp_byte_cnt_reg[7] (
	.clk(outclk_wire_0),
	.d(\Add4~25_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[7]~5_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(load_next_out_cmd1),
	.q(\out_uncomp_byte_cnt_reg[7]~q ),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[7] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[7] .power_up = "low";

cyclonev_lcell_comb \Add4~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\out_uncomp_byte_cnt_reg[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~26 ),
	.sharein(\Add4~27 ),
	.combout(),
	.sumout(\Add4~21_sumout ),
	.cout(),
	.shareout());
defparam \Add4~21 .extended_lut = "off";
defparam \Add4~21 .lut_mask = 64'h000000000000FF00;
defparam \Add4~21 .shared_arith = "on";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[8]~4 (
	.dataa(!WideOr0),
	.datab(!wrfull3),
	.datac(!wrfull2),
	.datad(!nxt_uncomp_subburst_byte_cnt),
	.datae(!\out_uncomp_byte_cnt_reg[8]~q ),
	.dataf(!\new_burst_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[8]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[8]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[8]~4 .lut_mask = 64'h005DFFFF0000FFA2;
defparam \nxt_uncomp_subburst_byte_cnt[8]~4 .shared_arith = "off";

dffeas \out_uncomp_byte_cnt_reg[8] (
	.clk(outclk_wire_0),
	.d(\Add4~21_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[8]~4_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(load_next_out_cmd1),
	.q(\out_uncomp_byte_cnt_reg[8]~q ),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[8] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[8] .power_up = "low";

cyclonev_lcell_comb \WideOr0~5 (
	.dataa(!\out_uncomp_byte_cnt_reg[8]~q ),
	.datab(!\out_uncomp_byte_cnt_reg[7]~q ),
	.datac(!\out_uncomp_byte_cnt_reg[2]~q ),
	.datad(!\out_uncomp_byte_cnt_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~5 .extended_lut = "off";
defparam \WideOr0~5 .lut_mask = 64'h8000800080008000;
defparam \WideOr0~5 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~1 (
	.dataa(!WideOr0),
	.datab(!wrfull3),
	.datac(!wrfull2),
	.datad(!nxt_uncomp_subburst_byte_cnt),
	.datae(!\new_burst_reg~q ),
	.dataf(!\WideOr0~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~1 .extended_lut = "off";
defparam \WideOr0~1 .lut_mask = 64'hFFFFFFA2005D0000;
defparam \WideOr0~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\Add4~1_sumout ),
	.datac(!\Add4~5_sumout ),
	.datad(!\Add4~9_sumout ),
	.datae(!\WideOr0~0_combout ),
	.dataf(!\WideOr0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~2 .extended_lut = "off";
defparam \WideOr0~2 .lut_mask = 64'hD555800080008000;
defparam \WideOr0~2 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\Add4~13_sumout ),
	.datac(!\Add4~17_sumout ),
	.datad(!\Add4~21_sumout ),
	.datae(!\Add4~25_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~3 .extended_lut = "off";
defparam \WideOr0~3 .lut_mask = 64'h2AAAAAAA2AAAAAAA;
defparam \WideOr0~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!nxt_in_ready),
	.datab(!\state.ST_IDLE~q ),
	.datac(!\in_valid~0_combout ),
	.datad(!in_eop_reg1),
	.datae(!\WideOr0~2_combout ),
	.dataf(!\WideOr0~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h0C0EAE0E0C0E0C0E;
defparam \Selector2~0 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(outclk_wire_0),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector3~1 (
	.dataa(!nxt_in_ready),
	.datab(!in_eop_reg1),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!\WideOr0~0_combout ),
	.datae(!\WideOr0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~1 .extended_lut = "off";
defparam \Selector3~1 .lut_mask = 64'h8088888880888888;
defparam \Selector3~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\Add4~1_sumout ),
	.datac(!\Add4~5_sumout ),
	.datad(!\Add4~9_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~2 .extended_lut = "off";
defparam \Selector3~2 .lut_mask = 64'h8000800080008000;
defparam \Selector3~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!\Add4~13_sumout ),
	.datab(!\Add4~17_sumout ),
	.datac(!\Add4~21_sumout ),
	.datad(!\Add4~25_sumout ),
	.datae(!\Selector3~1_combout ),
	.dataf(!\Selector3~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h0000FFFF00007FFF;
defparam \Selector3~0 .shared_arith = "off";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(outclk_wire_0),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\state.ST_UNCOMP_WR_SUBBURST~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready),
	.datac(!out_valid_reg1),
	.datad(!cp_ready),
	.datae(!mem_used_1),
	.dataf(!\in_valid~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h00000000D1DDD1D1;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_burstwrap[2]~0 (
	.dataa(!sink0_data[68]),
	.datab(!h2f_AWBURST_0),
	.datac(!h2f_AWBURST_1),
	.datad(!LessThan12),
	.datae(!Add4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_burstwrap[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_burstwrap[2]~0 .extended_lut = "off";
defparam \nxt_out_burstwrap[2]~0 .lut_mask = 64'h1511555115115551;
defparam \nxt_out_burstwrap[2]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(outclk_wire_0),
	.d(\nxt_out_burstwrap[2]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_out_burstwrap[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\in_burstwrap_reg[2]~q ),
	.datac(!\nxt_out_burstwrap[2]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_burstwrap[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_burstwrap[2]~1 .extended_lut = "off";
defparam \nxt_out_burstwrap[2]~1 .lut_mask = 64'h2727272727272727;
defparam \nxt_out_burstwrap[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!\d0_int_nxt_addr[2]~0_combout ),
	.datab(!\nxt_out_burstwrap[2]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h4444444444444444;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!in_data_reg_90),
	.datac(!in_data_reg_91),
	.datad(!sink0_data[91]),
	.datae(!sink0_data[90]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h085D0808085D0808;
defparam \ShiftLeft0~0 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!in_data_reg_90),
	.datac(!in_data_reg_91),
	.datad(!sink0_data[91]),
	.datae(!sink0_data[90]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h2020752020207520;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(outclk_wire_0),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_burstwrap[0]~5 (
	.dataa(!sink0_data[68]),
	.datab(!Selector8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_burstwrap[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_burstwrap[0]~5 .extended_lut = "off";
defparam \nxt_out_burstwrap[0]~5 .lut_mask = 64'h4444444444444444;
defparam \nxt_out_burstwrap[0]~5 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(outclk_wire_0),
	.d(\nxt_out_burstwrap[0]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_out_burstwrap[0]~6 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\in_burstwrap_reg[0]~q ),
	.datac(!\nxt_out_burstwrap[0]~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_burstwrap[0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_burstwrap[0]~6 .extended_lut = "off";
defparam \nxt_out_burstwrap[0]~6 .lut_mask = 64'h2727272727272727;
defparam \nxt_out_burstwrap[0]~6 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!\d0_int_nxt_addr[0]~3_combout ),
	.datab(!\nxt_out_burstwrap[0]~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h4444444444444444;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_data_36),
	.datac(!\Add0~13_sumout ),
	.datad(!\align_address_to_size|LessThan0~0_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'h0011AABB0A1BAABB;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[0]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_out_burstwrap[1]~4 (
	.dataa(!sink0_data[68]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!Selector7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_burstwrap[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_burstwrap[1]~4 .extended_lut = "off";
defparam \nxt_out_burstwrap[1]~4 .lut_mask = 64'h1D0C1D0C1D0C1D0C;
defparam \nxt_out_burstwrap[1]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!\d0_int_nxt_addr[1]~2_combout ),
	.datab(!\nxt_out_burstwrap[1]~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h4444444444444444;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \out_addr_reg~0 (
	.dataa(!\Add0~9_sumout ),
	.datab(!\int_nxt_addr_reg[1]~q ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_addr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_addr_reg~0 .extended_lut = "off";
defparam \out_addr_reg~0 .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \out_addr_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(gnd),
	.datac(!out_data_37),
	.datad(!sink0_data[91]),
	.datae(!\out_addr_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~2 .lut_mask = 64'hAFAA0500AFAA0500;
defparam \d0_int_nxt_addr[1]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!int_output_sel_0),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(!\in_burstwrap_reg[2]~q ),
	.datae(!\Add0~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~0 .lut_mask = 64'h1B1B1BBB1B1B1BBB;
defparam \d0_int_nxt_addr[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_burstwrap[3]~2 (
	.dataa(!sink0_data[68]),
	.datab(!h2f_AWBURST_0),
	.datac(!h2f_AWBURST_1),
	.datad(!Selector26),
	.datae(!Add41),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_burstwrap[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_burstwrap[3]~2 .extended_lut = "off";
defparam \nxt_out_burstwrap[3]~2 .lut_mask = 64'h1511555115115551;
defparam \nxt_out_burstwrap[3]~2 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(outclk_wire_0),
	.d(\nxt_out_burstwrap[3]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_out_burstwrap[3]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\in_burstwrap_reg[3]~q ),
	.datac(!\nxt_out_burstwrap[3]~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_burstwrap[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_burstwrap[3]~3 .extended_lut = "off";
defparam \nxt_out_burstwrap[3]~3 .lut_mask = 64'h2727272727272727;
defparam \nxt_out_burstwrap[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!\d0_int_nxt_addr[3]~1_combout ),
	.datab(!\nxt_out_burstwrap[3]~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h4444444444444444;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!in_data_reg_91),
	.datab(!in_data_reg_90),
	.datac(!\new_burst_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h1010101010101010;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(load_next_out_cmd1),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!int_output_sel_1),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(!\in_burstwrap_reg[3]~q ),
	.datae(!\Add0~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~1 .lut_mask = 64'h1B1B1BBB1B1B1BBB;
defparam \d0_int_nxt_addr[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_addr_reg~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_data_37),
	.datac(!\out_addr_reg~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_addr_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_addr_reg~1 .extended_lut = "off";
defparam \out_addr_reg~1 .lut_mask = 64'hB1B1B1B1B1B1B1B1;
defparam \out_addr_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \out_addr_reg~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_data_36),
	.datac(!\Add0~13_sumout ),
	.datad(!\int_nxt_addr_reg[0]~q ),
	.datae(!\in_burstwrap_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_addr_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_addr_reg~2 .extended_lut = "off";
defparam \out_addr_reg~2 .lut_mask = 64'h11BB1BBB11BB1BBB;
defparam \out_addr_reg~2 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_address_alignment_1 (
	new_burst_reg,
	in_data_reg_90,
	in_data_reg_91,
	out_data_90,
	out_data_91,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	in_data_reg_90;
input 	in_data_reg_91;
input 	out_data_90;
input 	out_data_91;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!in_data_reg_90),
	.datac(!in_data_reg_91),
	.datad(!out_data_91),
	.datae(!out_data_90),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hD5808080D5808080;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_burst_adapter_1 (
	outclk_wire_0,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_5,
	int_nxt_addr_reg_dly_6,
	int_nxt_addr_reg_dly_7,
	int_nxt_addr_reg_dly_8,
	int_nxt_addr_reg_dly_9,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_7,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_8,
	out_uncomp_byte_cnt_reg_5,
	out_burstwrap_reg_2,
	out_burstwrap_reg_3,
	out_addr_reg_1,
	out_burstwrap_reg_1,
	out_addr_reg_0,
	out_burstwrap_reg_0,
	Mux4,
	Mux5,
	Mux6,
	Mux7,
	Mux8,
	Mux9,
	Mux10,
	Mux11,
	Mux12,
	Mux13,
	Mux14,
	Mux15,
	Mux16,
	Mux17,
	Mux18,
	Mux19,
	Mux20,
	Mux21,
	Mux22,
	Mux23,
	Mux24,
	Mux25,
	Mux26,
	Mux27,
	Mux28,
	Mux29,
	Mux30,
	Mux31,
	Mux32,
	Mux33,
	Mux34,
	Mux35,
	in_ready_hold,
	saved_grant_1,
	saved_grant_0,
	src_data_198,
	src_data_199,
	src_data_200,
	stateST_COMP_TRANS,
	in_narrow_reg,
	always12,
	in_data_reg_91,
	in_data_reg_90,
	in_byteen_reg_2,
	source0_data_34,
	in_byteen_reg_0,
	source0_data_32,
	in_byteen_reg_1,
	source0_data_33,
	in_byteen_reg_3,
	source0_data_35,
	source0_data_351,
	mem_used_1,
	cp_ready,
	in_eop_reg,
	new_burst_reg,
	in_bytecount_reg_zero,
	nxt_in_ready,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	ShiftLeft1,
	source0_data_352,
	WideOr0,
	nxt_in_ready2,
	in_data_reg_68,
	in_data_reg_0,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	r_sync_rst,
	WideOr1,
	use_reg,
	nxt_out_eop,
	out_data_91,
	out_data_90,
	src_payload,
	src_data_190,
	out_data_37,
	src_payload1,
	src_data_189,
	out_data_36,
	int_output_sel_0,
	Mux1,
	Mux3,
	Mux2,
	Mux0,
	in_data_reg_69,
	cp_ready1,
	out_endofpacket,
	out_data_74,
	out_data_79,
	out_data_76,
	out_data_77,
	out_data_78,
	out_data_80,
	out_data_75,
	cp_ready2,
	out_byte_cnt_reg_2,
	src_valid,
	out_data_7,
	out_data_6,
	out_data_4,
	out_data_5,
	in_data_reg_122,
	in_data_reg_123,
	in_data_reg_124,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	in_data_reg_104,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	src_payload2,
	src_data_191,
	src_payload3,
	src_data_192,
	src_data_193,
	src_data_1931,
	address_reg_4,
	src_payload4,
	src_data_194,
	src_data_1941,
	address_reg_5,
	src_payload5,
	src_data_195,
	src_data_1951,
	address_reg_6,
	src_payload6,
	src_data_196,
	src_data_1961,
	address_reg_7,
	src_payload7,
	src_data_197,
	src_data_1971,
	out_data_44,
	out_data_45,
	src_data_1901,
	src_data_1891,
	src_data_209,
	src_data_210,
	src_data_211,
	src_data_212,
	src_data_213,
	src_data_214,
	src_data_215,
	src_data_216,
	src_data_217,
	src_data_218,
	src_data_219,
	src_data_220,
	src_data_1911,
	src_data_1921,
	src_data_1932,
	src_data_1942,
	src_data_1952,
	src_data_1962,
	src_data_1972,
	int_output_sel_1)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_5;
output 	int_nxt_addr_reg_dly_6;
output 	int_nxt_addr_reg_dly_7;
output 	int_nxt_addr_reg_dly_8;
output 	int_nxt_addr_reg_dly_9;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_7;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_8;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_burstwrap_reg_2;
output 	out_burstwrap_reg_3;
output 	out_addr_reg_1;
output 	out_burstwrap_reg_1;
output 	out_addr_reg_0;
output 	out_burstwrap_reg_0;
input 	Mux4;
input 	Mux5;
input 	Mux6;
input 	Mux7;
input 	Mux8;
input 	Mux9;
input 	Mux10;
input 	Mux11;
input 	Mux12;
input 	Mux13;
input 	Mux14;
input 	Mux15;
input 	Mux16;
input 	Mux17;
input 	Mux18;
input 	Mux19;
input 	Mux20;
input 	Mux21;
input 	Mux22;
input 	Mux23;
input 	Mux24;
input 	Mux25;
input 	Mux26;
input 	Mux27;
input 	Mux28;
input 	Mux29;
input 	Mux30;
input 	Mux31;
input 	Mux32;
input 	Mux33;
input 	Mux34;
input 	Mux35;
input 	in_ready_hold;
input 	saved_grant_1;
input 	saved_grant_0;
input 	src_data_198;
input 	src_data_199;
input 	src_data_200;
output 	stateST_COMP_TRANS;
output 	in_narrow_reg;
output 	always12;
output 	in_data_reg_91;
output 	in_data_reg_90;
output 	in_byteen_reg_2;
output 	source0_data_34;
output 	in_byteen_reg_0;
output 	source0_data_32;
output 	in_byteen_reg_1;
output 	source0_data_33;
output 	in_byteen_reg_3;
output 	source0_data_35;
output 	source0_data_351;
input 	mem_used_1;
input 	cp_ready;
output 	in_eop_reg;
output 	new_burst_reg;
output 	in_bytecount_reg_zero;
output 	nxt_in_ready;
output 	out_valid_reg;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
output 	ShiftLeft1;
output 	source0_data_352;
input 	WideOr0;
output 	nxt_in_ready2;
output 	in_data_reg_68;
output 	in_data_reg_0;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
input 	r_sync_rst;
input 	WideOr1;
input 	use_reg;
output 	nxt_out_eop;
input 	out_data_91;
input 	out_data_90;
input 	src_payload;
input 	src_data_190;
input 	out_data_37;
input 	src_payload1;
input 	src_data_189;
input 	out_data_36;
input 	int_output_sel_0;
input 	Mux1;
input 	Mux3;
input 	Mux2;
input 	Mux0;
output 	in_data_reg_69;
input 	cp_ready1;
input 	out_endofpacket;
input 	out_data_74;
input 	out_data_79;
input 	out_data_76;
input 	out_data_77;
input 	out_data_78;
input 	out_data_80;
input 	out_data_75;
input 	cp_ready2;
output 	out_byte_cnt_reg_2;
input 	src_valid;
input 	out_data_7;
input 	out_data_6;
input 	out_data_4;
input 	out_data_5;
output 	in_data_reg_122;
output 	in_data_reg_123;
output 	in_data_reg_124;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
output 	in_data_reg_104;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
input 	src_payload2;
input 	src_data_191;
input 	src_payload3;
input 	src_data_192;
input 	src_data_193;
input 	src_data_1931;
input 	address_reg_4;
input 	src_payload4;
input 	src_data_194;
input 	src_data_1941;
input 	address_reg_5;
input 	src_payload5;
input 	src_data_195;
input 	src_data_1951;
input 	address_reg_6;
input 	src_payload6;
input 	src_data_196;
input 	src_data_1961;
input 	address_reg_7;
input 	src_payload7;
input 	src_data_197;
input 	src_data_1971;
input 	out_data_44;
input 	out_data_45;
input 	src_data_1901;
input 	src_data_1891;
input 	src_data_209;
input 	src_data_210;
input 	src_data_211;
input 	src_data_212;
input 	src_data_213;
input 	src_data_214;
input 	src_data_215;
input 	src_data_216;
input 	src_data_217;
input 	src_data_218;
input 	src_data_219;
input 	src_data_220;
input 	src_data_1911;
input 	src_data_1921;
input 	src_data_1932;
input 	src_data_1942;
input 	src_data_1952;
input 	src_data_1962;
input 	src_data_1972;
input 	int_output_sel_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altera_merlin_burst_adapter_13_1_1 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.outclk_wire_0(outclk_wire_0),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_4(int_nxt_addr_reg_dly_4),
	.int_nxt_addr_reg_dly_5(int_nxt_addr_reg_dly_5),
	.int_nxt_addr_reg_dly_6(int_nxt_addr_reg_dly_6),
	.int_nxt_addr_reg_dly_7(int_nxt_addr_reg_dly_7),
	.int_nxt_addr_reg_dly_8(int_nxt_addr_reg_dly_8),
	.int_nxt_addr_reg_dly_9(int_nxt_addr_reg_dly_9),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_7(out_uncomp_byte_cnt_reg_7),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_8(out_uncomp_byte_cnt_reg_8),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_burstwrap_reg_2(out_burstwrap_reg_2),
	.out_burstwrap_reg_3(out_burstwrap_reg_3),
	.out_addr_reg_1(out_addr_reg_1),
	.out_burstwrap_reg_1(out_burstwrap_reg_1),
	.out_addr_reg_0(out_addr_reg_0),
	.out_burstwrap_reg_0(out_burstwrap_reg_0),
	.sink0_data({src_data_200,src_data_199,src_data_198,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_220,src_data_219,src_data_218,src_data_217,src_data_216,src_data_215,src_data_214,src_data_213,src_data_212,src_data_211,src_data_210,src_data_209,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,out_data_91,out_data_90,
src_data_1972,src_data_1962,src_data_1952,src_data_1942,src_data_1932,src_data_1921,src_data_1911,src_data_1901,src_data_1891,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,Mux0,Mux1,Mux2,Mux3,Mux4,Mux5,Mux6,Mux7,Mux8,Mux9,Mux10,Mux11,Mux12,Mux13,Mux14,Mux15,Mux16,Mux17,Mux18,Mux19,Mux20,Mux21,Mux22,Mux23,Mux24,Mux25,Mux26,Mux27,Mux28,Mux29,Mux30,Mux31,Mux32,Mux33,Mux34,Mux35}),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.in_narrow_reg1(in_narrow_reg),
	.always12(always12),
	.in_data_reg_91(in_data_reg_91),
	.in_data_reg_90(in_data_reg_90),
	.in_byteen_reg_2(in_byteen_reg_2),
	.source0_data_34(source0_data_34),
	.in_byteen_reg_0(in_byteen_reg_0),
	.source0_data_32(source0_data_32),
	.in_byteen_reg_1(in_byteen_reg_1),
	.source0_data_33(source0_data_33),
	.in_byteen_reg_3(in_byteen_reg_3),
	.source0_data_35(source0_data_35),
	.source0_data_351(source0_data_351),
	.mem_used_1(mem_used_1),
	.cp_ready(cp_ready),
	.in_eop_reg1(in_eop_reg),
	.new_burst_reg1(new_burst_reg),
	.in_bytecount_reg_zero1(in_bytecount_reg_zero),
	.nxt_in_ready(nxt_in_ready),
	.out_valid_reg1(out_valid_reg),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.ShiftLeft1(ShiftLeft1),
	.source0_data_352(source0_data_352),
	.WideOr0(WideOr0),
	.nxt_in_ready2(nxt_in_ready2),
	.in_data_reg_68(in_data_reg_68),
	.in_data_reg_0(in_data_reg_0),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_24(in_data_reg_24),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_31(in_data_reg_31),
	.r_sync_rst(r_sync_rst),
	.WideOr1(WideOr1),
	.use_reg(use_reg),
	.nxt_out_eop(nxt_out_eop),
	.src_payload(src_payload),
	.src_data_190(src_data_190),
	.out_data_37(out_data_37),
	.src_payload1(src_payload1),
	.src_data_189(src_data_189),
	.out_data_36(out_data_36),
	.int_output_sel_0(int_output_sel_0),
	.in_data_reg_69(in_data_reg_69),
	.cp_ready1(cp_ready1),
	.sink0_endofpacket(out_endofpacket),
	.out_data_74(out_data_74),
	.out_data_79(out_data_79),
	.out_data_76(out_data_76),
	.out_data_77(out_data_77),
	.out_data_78(out_data_78),
	.out_data_80(out_data_80),
	.out_data_75(out_data_75),
	.cp_ready2(cp_ready2),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.src_valid(src_valid),
	.out_data_7(out_data_7),
	.out_data_6(out_data_6),
	.out_data_4(out_data_4),
	.out_data_5(out_data_5),
	.in_data_reg_122(in_data_reg_122),
	.in_data_reg_123(in_data_reg_123),
	.in_data_reg_124(in_data_reg_124),
	.in_data_reg_101(in_data_reg_101),
	.in_data_reg_102(in_data_reg_102),
	.in_data_reg_103(in_data_reg_103),
	.in_data_reg_104(in_data_reg_104),
	.in_data_reg_105(in_data_reg_105),
	.in_data_reg_106(in_data_reg_106),
	.in_data_reg_107(in_data_reg_107),
	.in_data_reg_108(in_data_reg_108),
	.in_data_reg_109(in_data_reg_109),
	.in_data_reg_110(in_data_reg_110),
	.in_data_reg_111(in_data_reg_111),
	.in_data_reg_112(in_data_reg_112),
	.src_payload2(src_payload2),
	.src_data_191(src_data_191),
	.src_payload3(src_payload3),
	.src_data_192(src_data_192),
	.src_data_193(src_data_193),
	.src_data_1931(src_data_1931),
	.address_reg_4(address_reg_4),
	.src_payload4(src_payload4),
	.src_data_194(src_data_194),
	.src_data_1941(src_data_1941),
	.address_reg_5(address_reg_5),
	.src_payload5(src_payload5),
	.src_data_195(src_data_195),
	.src_data_1951(src_data_1951),
	.address_reg_6(address_reg_6),
	.src_payload6(src_payload6),
	.src_data_196(src_data_196),
	.src_data_1961(src_data_1961),
	.address_reg_7(address_reg_7),
	.src_payload7(src_payload7),
	.src_data_197(src_data_197),
	.src_data_1971(src_data_1971),
	.out_data_44(out_data_44),
	.out_data_45(out_data_45),
	.int_output_sel_1(int_output_sel_1));

endmodule

module Computer_System_altera_merlin_burst_adapter_13_1_1 (
	outclk_wire_0,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_5,
	int_nxt_addr_reg_dly_6,
	int_nxt_addr_reg_dly_7,
	int_nxt_addr_reg_dly_8,
	int_nxt_addr_reg_dly_9,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_7,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_8,
	out_uncomp_byte_cnt_reg_5,
	out_burstwrap_reg_2,
	out_burstwrap_reg_3,
	out_addr_reg_1,
	out_burstwrap_reg_1,
	out_addr_reg_0,
	out_burstwrap_reg_0,
	sink0_data,
	in_ready_hold,
	stateST_COMP_TRANS,
	in_narrow_reg1,
	always12,
	in_data_reg_91,
	in_data_reg_90,
	in_byteen_reg_2,
	source0_data_34,
	in_byteen_reg_0,
	source0_data_32,
	in_byteen_reg_1,
	source0_data_33,
	in_byteen_reg_3,
	source0_data_35,
	source0_data_351,
	mem_used_1,
	cp_ready,
	in_eop_reg1,
	new_burst_reg1,
	in_bytecount_reg_zero1,
	nxt_in_ready,
	out_valid_reg1,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	ShiftLeft1,
	source0_data_352,
	WideOr0,
	nxt_in_ready2,
	in_data_reg_68,
	in_data_reg_0,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	r_sync_rst,
	WideOr1,
	use_reg,
	nxt_out_eop,
	src_payload,
	src_data_190,
	out_data_37,
	src_payload1,
	src_data_189,
	out_data_36,
	int_output_sel_0,
	in_data_reg_69,
	cp_ready1,
	sink0_endofpacket,
	out_data_74,
	out_data_79,
	out_data_76,
	out_data_77,
	out_data_78,
	out_data_80,
	out_data_75,
	cp_ready2,
	out_byte_cnt_reg_2,
	src_valid,
	out_data_7,
	out_data_6,
	out_data_4,
	out_data_5,
	in_data_reg_122,
	in_data_reg_123,
	in_data_reg_124,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	in_data_reg_104,
	in_data_reg_105,
	in_data_reg_106,
	in_data_reg_107,
	in_data_reg_108,
	in_data_reg_109,
	in_data_reg_110,
	in_data_reg_111,
	in_data_reg_112,
	src_payload2,
	src_data_191,
	src_payload3,
	src_data_192,
	src_data_193,
	src_data_1931,
	address_reg_4,
	src_payload4,
	src_data_194,
	src_data_1941,
	address_reg_5,
	src_payload5,
	src_data_195,
	src_data_1951,
	address_reg_6,
	src_payload6,
	src_data_196,
	src_data_1961,
	address_reg_7,
	src_payload7,
	src_data_197,
	src_data_1971,
	out_data_44,
	out_data_45,
	int_output_sel_1)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_5;
output 	int_nxt_addr_reg_dly_6;
output 	int_nxt_addr_reg_dly_7;
output 	int_nxt_addr_reg_dly_8;
output 	int_nxt_addr_reg_dly_9;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_7;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_8;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_burstwrap_reg_2;
output 	out_burstwrap_reg_3;
output 	out_addr_reg_1;
output 	out_burstwrap_reg_1;
output 	out_addr_reg_0;
output 	out_burstwrap_reg_0;
input 	[124:0] sink0_data;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
output 	in_narrow_reg1;
output 	always12;
output 	in_data_reg_91;
output 	in_data_reg_90;
output 	in_byteen_reg_2;
output 	source0_data_34;
output 	in_byteen_reg_0;
output 	source0_data_32;
output 	in_byteen_reg_1;
output 	source0_data_33;
output 	in_byteen_reg_3;
output 	source0_data_35;
output 	source0_data_351;
input 	mem_used_1;
input 	cp_ready;
output 	in_eop_reg1;
output 	new_burst_reg1;
output 	in_bytecount_reg_zero1;
output 	nxt_in_ready;
output 	out_valid_reg1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
output 	ShiftLeft1;
output 	source0_data_352;
input 	WideOr0;
output 	nxt_in_ready2;
output 	in_data_reg_68;
output 	in_data_reg_0;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
input 	r_sync_rst;
input 	WideOr1;
input 	use_reg;
output 	nxt_out_eop;
input 	src_payload;
input 	src_data_190;
input 	out_data_37;
input 	src_payload1;
input 	src_data_189;
input 	out_data_36;
input 	int_output_sel_0;
output 	in_data_reg_69;
input 	cp_ready1;
input 	sink0_endofpacket;
input 	out_data_74;
input 	out_data_79;
input 	out_data_76;
input 	out_data_77;
input 	out_data_78;
input 	out_data_80;
input 	out_data_75;
input 	cp_ready2;
output 	out_byte_cnt_reg_2;
input 	src_valid;
input 	out_data_7;
input 	out_data_6;
input 	out_data_4;
input 	out_data_5;
output 	in_data_reg_122;
output 	in_data_reg_123;
output 	in_data_reg_124;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
output 	in_data_reg_104;
output 	in_data_reg_105;
output 	in_data_reg_106;
output 	in_data_reg_107;
output 	in_data_reg_108;
output 	in_data_reg_109;
output 	in_data_reg_110;
output 	in_data_reg_111;
output 	in_data_reg_112;
input 	src_payload2;
input 	src_data_191;
input 	src_payload3;
input 	src_data_192;
input 	src_data_193;
input 	src_data_1931;
input 	address_reg_4;
input 	src_payload4;
input 	src_data_194;
input 	src_data_1941;
input 	address_reg_5;
input 	src_payload5;
input 	src_data_195;
input 	src_data_1951;
input 	address_reg_6;
input 	src_payload6;
input 	src_data_196;
input 	src_data_1961;
input 	address_reg_7;
input 	src_payload7;
input 	src_data_197;
input 	src_data_1971;
input 	out_data_44;
input 	out_data_45;
input 	int_output_sel_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|out_data[1]~combout ;
wire \align_address_to_size|LessThan0~0_combout ;
wire \align_address_to_size|out_data[0]~combout ;
wire \ShiftLeft0~1_combout ;
wire \load_next_out_cmd~combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~5_sumout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~1_combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \int_nxt_addr_with_offset[0]~combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~0_combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \int_nxt_addr_with_offset[1]~combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~2 ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~2_combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \int_nxt_addr_with_offset[2]~combout ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~3_combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \int_nxt_addr_with_offset[3]~combout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \in_burstwrap_reg[4]~q ;
wire \d0_int_nxt_addr[4]~0_combout ;
wire \nxt_addr[4]~4_combout ;
wire \int_nxt_addr_reg[4]~q ;
wire \int_nxt_addr_with_offset[4]~combout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \in_burstwrap_reg[5]~q ;
wire \d0_int_nxt_addr[5]~1_combout ;
wire \nxt_addr[5]~5_combout ;
wire \int_nxt_addr_reg[5]~q ;
wire \int_nxt_addr_with_offset[5]~combout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \in_burstwrap_reg[6]~q ;
wire \d0_int_nxt_addr[6]~2_combout ;
wire \nxt_addr[6]~6_combout ;
wire \int_nxt_addr_reg[6]~q ;
wire \int_nxt_addr_with_offset[6]~combout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \in_burstwrap_reg[7]~q ;
wire \d0_int_nxt_addr[7]~3_combout ;
wire \nxt_addr[7]~7_combout ;
wire \int_nxt_addr_reg[7]~q ;
wire \int_nxt_addr_with_offset[7]~combout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \in_burstwrap_reg[8]~q ;
wire \nxt_addr[8]~8_combout ;
wire \int_nxt_addr_reg[8]~q ;
wire \int_nxt_addr_with_offset[8]~combout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \nxt_addr[9]~9_combout ;
wire \int_nxt_addr_reg[9]~q ;
wire \int_nxt_addr_with_offset[9]~combout ;
wire \Add4~6 ;
wire \Add4~7 ;
wire \Add4~10 ;
wire \Add4~11 ;
wire \Add4~14 ;
wire \Add4~15 ;
wire \Add4~18 ;
wire \Add4~19 ;
wire \Add4~21_sumout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[7]~3_combout ;
wire \WideOr0~0_combout ;
wire \WideOr0~1_combout ;
wire \Add4~22 ;
wire \Add4~23 ;
wire \Add4~26 ;
wire \Add4~27 ;
wire \Add4~1_sumout ;
wire \Add4~5_sumout ;
wire \Add4~9_sumout ;
wire \Add4~13_sumout ;
wire \Add4~17_sumout ;
wire \Add4~25_sumout ;
wire \WideOr0~2_combout ;
wire \nxt_in_ready~1_combout ;
wire \Selector3~0_combout ;
wire \nxt_out_eop~0_combout ;
wire \Selector0~0_combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \Selector2~3_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \nxt_uncomp_subburst_byte_cnt[4]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[8]~5_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~6_combout ;
wire \always10~0_combout ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \in_narrow_reg~0_combout ;
wire \new_burst_reg~0_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \Add1~17_sumout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \Add1~18 ;
wire \Add1~19 ;
wire \Add1~21_sumout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~22 ;
wire \Add1~23 ;
wire \Add1~25_sumout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~26 ;
wire \Add1~27 ;
wire \Add1~1_sumout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \Add1~2 ;
wire \Add1~3 ;
wire \Add1~5_sumout ;
wire \int_bytes_remaining_reg[7]~q ;
wire \Add1~6 ;
wire \Add1~7 ;
wire \Add1~9_sumout ;
wire \int_bytes_remaining_reg[8]~q ;
wire \Add1~10 ;
wire \Add1~11 ;
wire \Add1~13_sumout ;
wire \new_burst_reg~1_combout ;
wire \new_burst_reg~2_combout ;
wire \new_burst_reg~3_combout ;
wire \WideNor0~combout ;
wire \nxt_out_valid~0_combout ;
wire \WideOr0~3_combout ;
wire \Selector3~1_combout ;
wire \nxt_in_ready~3_combout ;


Computer_System_altera_merlin_address_alignment_2 align_address_to_size(
	.src_data_198(sink0_data[122]),
	.src_data_199(sink0_data[123]),
	.src_data_200(sink0_data[124]),
	.in_data_reg_91(in_data_reg_91),
	.in_data_reg_90(in_data_reg_90),
	.new_burst_reg(new_burst_reg1),
	.out_data_91(sink0_data[91]),
	.out_data_37(out_data_37),
	.out_data_1(\align_address_to_size|out_data[1]~combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ),
	.out_data_36(out_data_36),
	.out_data_0(\align_address_to_size|out_data[0]~combout ));

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(outclk_wire_0),
	.d(\int_nxt_addr_with_offset[2]~combout ),
	.asdata(int_output_sel_0),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(outclk_wire_0),
	.d(\int_nxt_addr_with_offset[3]~combout ),
	.asdata(int_output_sel_1),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[4] (
	.clk(outclk_wire_0),
	.d(\int_nxt_addr_with_offset[4]~combout ),
	.asdata(\d0_int_nxt_addr[4]~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_4),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[4] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[4] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[5] (
	.clk(outclk_wire_0),
	.d(\int_nxt_addr_with_offset[5]~combout ),
	.asdata(\d0_int_nxt_addr[5]~1_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_5),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[5] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[5] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[6] (
	.clk(outclk_wire_0),
	.d(\int_nxt_addr_with_offset[6]~combout ),
	.asdata(\d0_int_nxt_addr[6]~2_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_6),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[6] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[6] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[7] (
	.clk(outclk_wire_0),
	.d(\int_nxt_addr_with_offset[7]~combout ),
	.asdata(\d0_int_nxt_addr[7]~3_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_7),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[7] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[7] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[8] (
	.clk(outclk_wire_0),
	.d(\int_nxt_addr_with_offset[8]~combout ),
	.asdata(out_data_44),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_8),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[8] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[8] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[9] (
	.clk(outclk_wire_0),
	.d(\int_nxt_addr_with_offset[9]~combout ),
	.asdata(out_data_45),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_9),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[9] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[9] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(outclk_wire_0),
	.d(\Add4~21_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[6]~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(outclk_wire_0),
	.d(\Add4~5_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[2]~1_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(outclk_wire_0),
	.d(\Add4~9_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[7] (
	.clk(outclk_wire_0),
	.d(\Add4~25_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[7]~3_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_7),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[7] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[7] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(outclk_wire_0),
	.d(\Add4~13_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[8] (
	.clk(outclk_wire_0),
	.d(\Add4~1_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[8]~5_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_8),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[8] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[8] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(outclk_wire_0),
	.d(\Add4~17_sumout ),
	.asdata(\nxt_uncomp_subburst_byte_cnt[5]~6_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.ST_UNCOMP_TRANS~q ),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_burstwrap_reg[2] (
	.clk(outclk_wire_0),
	.d(\in_burstwrap_reg[2]~q ),
	.asdata(sink0_data[83]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\always10~0_combout ),
	.q(out_burstwrap_reg_2),
	.prn(vcc));
defparam \out_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \out_burstwrap_reg[2] .power_up = "low";

dffeas \out_burstwrap_reg[3] (
	.clk(outclk_wire_0),
	.d(\in_burstwrap_reg[3]~q ),
	.asdata(sink0_data[84]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\always10~0_combout ),
	.q(out_burstwrap_reg_3),
	.prn(vcc));
defparam \out_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \out_burstwrap_reg[3] .power_up = "low";

dffeas \out_addr_reg[1] (
	.clk(outclk_wire_0),
	.d(\int_nxt_addr_with_offset[1]~combout ),
	.asdata(out_data_37),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(out_addr_reg_1),
	.prn(vcc));
defparam \out_addr_reg[1] .is_wysiwyg = "true";
defparam \out_addr_reg[1] .power_up = "low";

dffeas \out_burstwrap_reg[1] (
	.clk(outclk_wire_0),
	.d(\in_burstwrap_reg[1]~q ),
	.asdata(sink0_data[82]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\always10~0_combout ),
	.q(out_burstwrap_reg_1),
	.prn(vcc));
defparam \out_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \out_burstwrap_reg[1] .power_up = "low";

dffeas \out_addr_reg[0] (
	.clk(outclk_wire_0),
	.d(\int_nxt_addr_with_offset[0]~combout ),
	.asdata(out_data_36),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(out_addr_reg_0),
	.prn(vcc));
defparam \out_addr_reg[0] .is_wysiwyg = "true";
defparam \out_addr_reg[0] .power_up = "low";

dffeas \out_burstwrap_reg[0] (
	.clk(outclk_wire_0),
	.d(\in_burstwrap_reg[0]~q ),
	.asdata(sink0_data[81]),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\always10~0_combout ),
	.q(out_burstwrap_reg_0),
	.prn(vcc));
defparam \out_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \out_burstwrap_reg[0] .power_up = "low";

dffeas \state.ST_COMP_TRANS (
	.clk(outclk_wire_0),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas in_narrow_reg(
	.clk(outclk_wire_0),
	.d(\in_narrow_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

cyclonev_lcell_comb \always12~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always12),
	.sumout(),
	.cout(),
	.shareout());
defparam \always12~0 .extended_lut = "off";
defparam \always12~0 .lut_mask = 64'h1111111111111111;
defparam \always12~0 .shared_arith = "off";

dffeas \in_data_reg[91] (
	.clk(outclk_wire_0),
	.d(sink0_data[91]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_91),
	.prn(vcc));
defparam \in_data_reg[91] .is_wysiwyg = "true";
defparam \in_data_reg[91] .power_up = "low";

dffeas \in_data_reg[90] (
	.clk(outclk_wire_0),
	.d(sink0_data[90]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_90),
	.prn(vcc));
defparam \in_data_reg[90] .is_wysiwyg = "true";
defparam \in_data_reg[90] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

cyclonev_lcell_comb \source0_data[34]~0 (
	.dataa(!always12),
	.datab(!in_data_reg_91),
	.datac(!in_data_reg_90),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(!\int_nxt_addr_reg_dly[0]~q ),
	.dataf(!in_byteen_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[34]~0 .extended_lut = "off";
defparam \source0_data[34]~0 .lut_mask = 64'h11551500BBFFBFAA;
defparam \source0_data[34]~0 .shared_arith = "off";

dffeas \in_byteen_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

cyclonev_lcell_comb \source0_data[32]~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg1),
	.datac(!\int_nxt_addr_reg_dly[1]~q ),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(!in_byteen_reg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[32]~1 .extended_lut = "off";
defparam \source0_data[32]~1 .lut_mask = 64'h1000FEEE1000FEEE;
defparam \source0_data[32]~1 .shared_arith = "off";

dffeas \in_byteen_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

cyclonev_lcell_comb \source0_data[33]~2 (
	.dataa(!always12),
	.datab(!in_data_reg_91),
	.datac(!in_data_reg_90),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(!\int_nxt_addr_reg_dly[0]~q ),
	.dataf(!in_byteen_reg_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[33]~2 .extended_lut = "off";
defparam \source0_data[33]~2 .lut_mask = 64'h15005500BFAAFFAA;
defparam \source0_data[33]~2 .shared_arith = "off";

dffeas \in_byteen_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

cyclonev_lcell_comb \source0_data[35]~3 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg1),
	.datac(!in_data_reg_91),
	.datad(!in_byteen_reg_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[35]~3 .extended_lut = "off";
defparam \source0_data[35]~3 .lut_mask = 64'h01EF01EF01EF01EF;
defparam \source0_data[35]~3 .shared_arith = "off";

cyclonev_lcell_comb \source0_data[35]~4 (
	.dataa(!always12),
	.datab(!in_data_reg_90),
	.datac(!\int_nxt_addr_reg_dly[1]~q ),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(!source0_data_35),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_351),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[35]~4 .extended_lut = "off";
defparam \source0_data[35]~4 .lut_mask = 64'h0105FFFF0105FFFF;
defparam \source0_data[35]~4 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(outclk_wire_0),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_eop_reg1),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

dffeas new_burst_reg(
	.clk(outclk_wire_0),
	.d(\new_burst_reg~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(new_burst_reg1),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

dffeas in_bytecount_reg_zero(
	.clk(outclk_wire_0),
	.d(\WideNor0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_bytecount_reg_zero1),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!cp_ready),
	.datac(gnd),
	.datad(!new_burst_reg1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h0011001100110011;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(outclk_wire_0),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(outclk_wire_0),
	.d(\Selector3~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~2 (
	.dataa(!in_ready_hold),
	.datab(!out_valid_reg1),
	.datac(!stateST_COMP_TRANS),
	.datad(!cp_ready),
	.datae(!\nxt_in_ready~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~2 .extended_lut = "off";
defparam \nxt_in_ready~2 .lut_mask = 64'h3303A3A33303A3A3;
defparam \nxt_in_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft1~0 (
	.dataa(!in_data_reg_91),
	.datab(!in_data_reg_90),
	.datac(!\int_nxt_addr_reg_dly[1]~q ),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft1),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft1~0 .extended_lut = "off";
defparam \ShiftLeft1~0 .lut_mask = 64'hA08FA08FA08FA08F;
defparam \ShiftLeft1~0 .shared_arith = "off";

cyclonev_lcell_comb \source0_data[35]~5 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg1),
	.datac(!in_data_reg_90),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(!\int_nxt_addr_reg_dly[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source0_data_352),
	.sumout(),
	.cout(),
	.shareout());
defparam \source0_data[35]~5 .extended_lut = "off";
defparam \source0_data[35]~5 .lut_mask = 64'h0001001100010011;
defparam \source0_data[35]~5 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~4 (
	.dataa(!out_valid_reg1),
	.datab(!stateST_COMP_TRANS),
	.datac(!cp_ready),
	.datad(gnd),
	.datae(!\nxt_out_eop~0_combout ),
	.dataf(!\nxt_in_ready~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~4 .extended_lut = "off";
defparam \nxt_in_ready~4 .lut_mask = 64'h11111010DDDDDCDC;
defparam \nxt_in_ready~4 .shared_arith = "off";

dffeas \in_data_reg[68] (
	.clk(outclk_wire_0),
	.d(sink0_data[68]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_68),
	.prn(vcc));
defparam \in_data_reg[68] .is_wysiwyg = "true";
defparam \in_data_reg[68] .power_up = "low";

dffeas \in_data_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \in_data_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_1),
	.prn(vcc));
defparam \in_data_reg[1] .is_wysiwyg = "true";
defparam \in_data_reg[1] .power_up = "low";

dffeas \in_data_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_2),
	.prn(vcc));
defparam \in_data_reg[2] .is_wysiwyg = "true";
defparam \in_data_reg[2] .power_up = "low";

dffeas \in_data_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_3),
	.prn(vcc));
defparam \in_data_reg[3] .is_wysiwyg = "true";
defparam \in_data_reg[3] .power_up = "low";

dffeas \in_data_reg[4] (
	.clk(outclk_wire_0),
	.d(sink0_data[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_4),
	.prn(vcc));
defparam \in_data_reg[4] .is_wysiwyg = "true";
defparam \in_data_reg[4] .power_up = "low";

dffeas \in_data_reg[5] (
	.clk(outclk_wire_0),
	.d(sink0_data[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_5),
	.prn(vcc));
defparam \in_data_reg[5] .is_wysiwyg = "true";
defparam \in_data_reg[5] .power_up = "low";

dffeas \in_data_reg[6] (
	.clk(outclk_wire_0),
	.d(sink0_data[6]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_6),
	.prn(vcc));
defparam \in_data_reg[6] .is_wysiwyg = "true";
defparam \in_data_reg[6] .power_up = "low";

dffeas \in_data_reg[7] (
	.clk(outclk_wire_0),
	.d(sink0_data[7]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_7),
	.prn(vcc));
defparam \in_data_reg[7] .is_wysiwyg = "true";
defparam \in_data_reg[7] .power_up = "low";

dffeas \in_data_reg[8] (
	.clk(outclk_wire_0),
	.d(sink0_data[8]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_8),
	.prn(vcc));
defparam \in_data_reg[8] .is_wysiwyg = "true";
defparam \in_data_reg[8] .power_up = "low";

dffeas \in_data_reg[9] (
	.clk(outclk_wire_0),
	.d(sink0_data[9]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_9),
	.prn(vcc));
defparam \in_data_reg[9] .is_wysiwyg = "true";
defparam \in_data_reg[9] .power_up = "low";

dffeas \in_data_reg[10] (
	.clk(outclk_wire_0),
	.d(sink0_data[10]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_10),
	.prn(vcc));
defparam \in_data_reg[10] .is_wysiwyg = "true";
defparam \in_data_reg[10] .power_up = "low";

dffeas \in_data_reg[11] (
	.clk(outclk_wire_0),
	.d(sink0_data[11]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_11),
	.prn(vcc));
defparam \in_data_reg[11] .is_wysiwyg = "true";
defparam \in_data_reg[11] .power_up = "low";

dffeas \in_data_reg[12] (
	.clk(outclk_wire_0),
	.d(sink0_data[12]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_12),
	.prn(vcc));
defparam \in_data_reg[12] .is_wysiwyg = "true";
defparam \in_data_reg[12] .power_up = "low";

dffeas \in_data_reg[13] (
	.clk(outclk_wire_0),
	.d(sink0_data[13]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_13),
	.prn(vcc));
defparam \in_data_reg[13] .is_wysiwyg = "true";
defparam \in_data_reg[13] .power_up = "low";

dffeas \in_data_reg[14] (
	.clk(outclk_wire_0),
	.d(sink0_data[14]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_14),
	.prn(vcc));
defparam \in_data_reg[14] .is_wysiwyg = "true";
defparam \in_data_reg[14] .power_up = "low";

dffeas \in_data_reg[15] (
	.clk(outclk_wire_0),
	.d(sink0_data[15]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_15),
	.prn(vcc));
defparam \in_data_reg[15] .is_wysiwyg = "true";
defparam \in_data_reg[15] .power_up = "low";

dffeas \in_data_reg[16] (
	.clk(outclk_wire_0),
	.d(sink0_data[16]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_16),
	.prn(vcc));
defparam \in_data_reg[16] .is_wysiwyg = "true";
defparam \in_data_reg[16] .power_up = "low";

dffeas \in_data_reg[17] (
	.clk(outclk_wire_0),
	.d(sink0_data[17]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_17),
	.prn(vcc));
defparam \in_data_reg[17] .is_wysiwyg = "true";
defparam \in_data_reg[17] .power_up = "low";

dffeas \in_data_reg[18] (
	.clk(outclk_wire_0),
	.d(sink0_data[18]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_18),
	.prn(vcc));
defparam \in_data_reg[18] .is_wysiwyg = "true";
defparam \in_data_reg[18] .power_up = "low";

dffeas \in_data_reg[19] (
	.clk(outclk_wire_0),
	.d(sink0_data[19]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_19),
	.prn(vcc));
defparam \in_data_reg[19] .is_wysiwyg = "true";
defparam \in_data_reg[19] .power_up = "low";

dffeas \in_data_reg[20] (
	.clk(outclk_wire_0),
	.d(sink0_data[20]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_20),
	.prn(vcc));
defparam \in_data_reg[20] .is_wysiwyg = "true";
defparam \in_data_reg[20] .power_up = "low";

dffeas \in_data_reg[21] (
	.clk(outclk_wire_0),
	.d(sink0_data[21]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_21),
	.prn(vcc));
defparam \in_data_reg[21] .is_wysiwyg = "true";
defparam \in_data_reg[21] .power_up = "low";

dffeas \in_data_reg[22] (
	.clk(outclk_wire_0),
	.d(sink0_data[22]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_22),
	.prn(vcc));
defparam \in_data_reg[22] .is_wysiwyg = "true";
defparam \in_data_reg[22] .power_up = "low";

dffeas \in_data_reg[23] (
	.clk(outclk_wire_0),
	.d(sink0_data[23]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_23),
	.prn(vcc));
defparam \in_data_reg[23] .is_wysiwyg = "true";
defparam \in_data_reg[23] .power_up = "low";

dffeas \in_data_reg[24] (
	.clk(outclk_wire_0),
	.d(sink0_data[24]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_24),
	.prn(vcc));
defparam \in_data_reg[24] .is_wysiwyg = "true";
defparam \in_data_reg[24] .power_up = "low";

dffeas \in_data_reg[25] (
	.clk(outclk_wire_0),
	.d(sink0_data[25]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_25),
	.prn(vcc));
defparam \in_data_reg[25] .is_wysiwyg = "true";
defparam \in_data_reg[25] .power_up = "low";

dffeas \in_data_reg[26] (
	.clk(outclk_wire_0),
	.d(sink0_data[26]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_26),
	.prn(vcc));
defparam \in_data_reg[26] .is_wysiwyg = "true";
defparam \in_data_reg[26] .power_up = "low";

dffeas \in_data_reg[27] (
	.clk(outclk_wire_0),
	.d(sink0_data[27]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_27),
	.prn(vcc));
defparam \in_data_reg[27] .is_wysiwyg = "true";
defparam \in_data_reg[27] .power_up = "low";

dffeas \in_data_reg[28] (
	.clk(outclk_wire_0),
	.d(sink0_data[28]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_28),
	.prn(vcc));
defparam \in_data_reg[28] .is_wysiwyg = "true";
defparam \in_data_reg[28] .power_up = "low";

dffeas \in_data_reg[29] (
	.clk(outclk_wire_0),
	.d(sink0_data[29]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_29),
	.prn(vcc));
defparam \in_data_reg[29] .is_wysiwyg = "true";
defparam \in_data_reg[29] .power_up = "low";

dffeas \in_data_reg[30] (
	.clk(outclk_wire_0),
	.d(sink0_data[30]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_30),
	.prn(vcc));
defparam \in_data_reg[30] .is_wysiwyg = "true";
defparam \in_data_reg[30] .power_up = "low";

dffeas \in_data_reg[31] (
	.clk(outclk_wire_0),
	.d(sink0_data[31]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_31),
	.prn(vcc));
defparam \in_data_reg[31] .is_wysiwyg = "true";
defparam \in_data_reg[31] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!cp_ready),
	.datac(!in_eop_reg1),
	.datad(!new_burst_reg1),
	.datae(!in_bytecount_reg_zero1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~1 .extended_lut = "off";
defparam \nxt_out_eop~1 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \nxt_out_eop~1 .shared_arith = "off";

dffeas \in_data_reg[69] (
	.clk(outclk_wire_0),
	.d(sink0_data[69]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_69),
	.prn(vcc));
defparam \in_data_reg[69] .is_wysiwyg = "true";
defparam \in_data_reg[69] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(outclk_wire_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \in_data_reg[122] (
	.clk(outclk_wire_0),
	.d(sink0_data[122]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_122),
	.prn(vcc));
defparam \in_data_reg[122] .is_wysiwyg = "true";
defparam \in_data_reg[122] .power_up = "low";

dffeas \in_data_reg[123] (
	.clk(outclk_wire_0),
	.d(sink0_data[123]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_123),
	.prn(vcc));
defparam \in_data_reg[123] .is_wysiwyg = "true";
defparam \in_data_reg[123] .power_up = "low";

dffeas \in_data_reg[124] (
	.clk(outclk_wire_0),
	.d(sink0_data[124]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_124),
	.prn(vcc));
defparam \in_data_reg[124] .is_wysiwyg = "true";
defparam \in_data_reg[124] .power_up = "low";

dffeas \in_data_reg[101] (
	.clk(outclk_wire_0),
	.d(sink0_data[101]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_101),
	.prn(vcc));
defparam \in_data_reg[101] .is_wysiwyg = "true";
defparam \in_data_reg[101] .power_up = "low";

dffeas \in_data_reg[102] (
	.clk(outclk_wire_0),
	.d(sink0_data[102]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_102),
	.prn(vcc));
defparam \in_data_reg[102] .is_wysiwyg = "true";
defparam \in_data_reg[102] .power_up = "low";

dffeas \in_data_reg[103] (
	.clk(outclk_wire_0),
	.d(sink0_data[103]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_103),
	.prn(vcc));
defparam \in_data_reg[103] .is_wysiwyg = "true";
defparam \in_data_reg[103] .power_up = "low";

dffeas \in_data_reg[104] (
	.clk(outclk_wire_0),
	.d(sink0_data[104]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_104),
	.prn(vcc));
defparam \in_data_reg[104] .is_wysiwyg = "true";
defparam \in_data_reg[104] .power_up = "low";

dffeas \in_data_reg[105] (
	.clk(outclk_wire_0),
	.d(sink0_data[105]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_105),
	.prn(vcc));
defparam \in_data_reg[105] .is_wysiwyg = "true";
defparam \in_data_reg[105] .power_up = "low";

dffeas \in_data_reg[106] (
	.clk(outclk_wire_0),
	.d(sink0_data[106]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_106),
	.prn(vcc));
defparam \in_data_reg[106] .is_wysiwyg = "true";
defparam \in_data_reg[106] .power_up = "low";

dffeas \in_data_reg[107] (
	.clk(outclk_wire_0),
	.d(sink0_data[107]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_107),
	.prn(vcc));
defparam \in_data_reg[107] .is_wysiwyg = "true";
defparam \in_data_reg[107] .power_up = "low";

dffeas \in_data_reg[108] (
	.clk(outclk_wire_0),
	.d(sink0_data[108]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_108),
	.prn(vcc));
defparam \in_data_reg[108] .is_wysiwyg = "true";
defparam \in_data_reg[108] .power_up = "low";

dffeas \in_data_reg[109] (
	.clk(outclk_wire_0),
	.d(sink0_data[109]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_109),
	.prn(vcc));
defparam \in_data_reg[109] .is_wysiwyg = "true";
defparam \in_data_reg[109] .power_up = "low";

dffeas \in_data_reg[110] (
	.clk(outclk_wire_0),
	.d(sink0_data[110]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_110),
	.prn(vcc));
defparam \in_data_reg[110] .is_wysiwyg = "true";
defparam \in_data_reg[110] .power_up = "low";

dffeas \in_data_reg[111] (
	.clk(outclk_wire_0),
	.d(sink0_data[111]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_111),
	.prn(vcc));
defparam \in_data_reg[111] .is_wysiwyg = "true";
defparam \in_data_reg[111] .power_up = "low";

dffeas \in_data_reg[112] (
	.clk(outclk_wire_0),
	.d(sink0_data[112]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_112),
	.prn(vcc));
defparam \in_data_reg[112] .is_wysiwyg = "true";
defparam \in_data_reg[112] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!in_data_reg_91),
	.datab(!in_data_reg_90),
	.datac(!new_burst_reg1),
	.datad(!sink0_data[91]),
	.datae(!sink0_data[90]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h404F4040404F4040;
defparam \ShiftLeft0~1 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!in_ready_hold),
	.datab(!out_valid_reg1),
	.datac(!source0_data_33),
	.datad(!WideOr0),
	.datae(!mem_used_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hDDFDCCCCDDFDCCCC;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!in_data_reg_91),
	.datab(!in_data_reg_90),
	.datac(!new_burst_reg1),
	.datad(!sink0_data[91]),
	.datae(!sink0_data[90]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h20202F2020202F20;
defparam \ShiftLeft0~0 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(outclk_wire_0),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready),
	.datac(!nxt_in_ready1),
	.datad(!WideOr1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0051005100510051;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[81]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0]~1 (
	.dataa(!new_burst_reg1),
	.datab(!sink0_data[81]),
	.datac(!\in_burstwrap_reg[0]~q ),
	.datad(!\int_nxt_addr_with_offset[0]~combout ),
	.datae(!\align_address_to_size|out_data[0]~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0]~1 .extended_lut = "off";
defparam \nxt_addr[0]~1 .lut_mask = 64'h00A044E400A044E4;
defparam \nxt_addr[0]~1 .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[0] (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~5_sumout ),
	.datac(!src_payload1),
	.datad(!src_data_189),
	.datae(!\in_burstwrap_reg[0]~q ),
	.dataf(!\int_nxt_addr_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[0] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[0] .lut_mask = 64'h01112333FFFFFFFF;
defparam \int_nxt_addr_with_offset[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(outclk_wire_0),
	.d(\int_nxt_addr_with_offset[0]~combout ),
	.asdata(\align_address_to_size|out_data[0]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[82]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1]~0 (
	.dataa(!new_burst_reg1),
	.datab(!sink0_data[82]),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\int_nxt_addr_with_offset[1]~combout ),
	.datae(!\align_address_to_size|out_data[1]~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1]~0 .extended_lut = "off";
defparam \nxt_addr[1]~0 .lut_mask = 64'h00A044E400A044E4;
defparam \nxt_addr[1]~0 .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[1] (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~1_sumout ),
	.datac(!src_payload),
	.datad(!src_data_190),
	.datae(!\in_burstwrap_reg[1]~q ),
	.dataf(!\int_nxt_addr_reg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[1] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[1] .lut_mask = 64'h01112333FFFFFFFF;
defparam \int_nxt_addr_with_offset[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(outclk_wire_0),
	.d(\int_nxt_addr_with_offset[1]~combout ),
	.asdata(\align_address_to_size|out_data[1]~combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[83]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2]~2 (
	.dataa(!new_burst_reg1),
	.datab(!int_output_sel_0),
	.datac(!sink0_data[83]),
	.datad(!\in_burstwrap_reg[2]~q ),
	.datae(!\int_nxt_addr_with_offset[2]~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2]~2 .extended_lut = "off";
defparam \nxt_addr[2]~2 .lut_mask = 64'h1010BA101010BA10;
defparam \nxt_addr[2]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[2] (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~9_sumout ),
	.datac(!src_payload2),
	.datad(!src_data_191),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\int_nxt_addr_reg[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[2] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[2] .lut_mask = 64'h01112333FFFFFFFF;
defparam \int_nxt_addr_with_offset[2] .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!new_burst_reg1),
	.datab(!in_data_reg_90),
	.datac(!in_data_reg_91),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h0202020202020202;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[84]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3]~3 (
	.dataa(!new_burst_reg1),
	.datab(!int_output_sel_1),
	.datac(!sink0_data[84]),
	.datad(!\in_burstwrap_reg[3]~q ),
	.datae(!\int_nxt_addr_with_offset[3]~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3]~3 .extended_lut = "off";
defparam \nxt_addr[3]~3 .lut_mask = 64'h1010BA101010BA10;
defparam \nxt_addr[3]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[3] (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~13_sumout ),
	.datac(!src_payload3),
	.datad(!src_data_192),
	.datae(!\in_burstwrap_reg[3]~q ),
	.dataf(!\int_nxt_addr_reg[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[3] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[3] .lut_mask = 64'h01112333FFFFFFFF;
defparam \int_nxt_addr_with_offset[3] .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \in_burstwrap_reg[4] (
	.clk(outclk_wire_0),
	.d(sink0_data[85]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[4]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[4] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[4] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[4]~0 (
	.dataa(!sink0_data[68]),
	.datab(!out_data_4),
	.datac(!use_reg),
	.datad(!address_reg_4),
	.datae(!src_payload4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[4]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[4]~0 .lut_mask = 64'h101FF0FF101FF0FF;
defparam \d0_int_nxt_addr[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[4]~4 (
	.dataa(!new_burst_reg1),
	.datab(!sink0_data[85]),
	.datac(!\in_burstwrap_reg[4]~q ),
	.datad(!\int_nxt_addr_with_offset[4]~combout ),
	.datae(!\d0_int_nxt_addr[4]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[4]~4 .extended_lut = "off";
defparam \nxt_addr[4]~4 .lut_mask = 64'h00A044E400A044E4;
defparam \nxt_addr[4]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg[4] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[4]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[4] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[4] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[4] (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~17_sumout ),
	.datac(!src_data_193),
	.datad(!src_data_1931),
	.datae(!\in_burstwrap_reg[4]~q ),
	.dataf(!\int_nxt_addr_reg[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[4] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[4] .lut_mask = 64'h01112333FFFFFFFF;
defparam \int_nxt_addr_with_offset[4] .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \in_burstwrap_reg[5] (
	.clk(outclk_wire_0),
	.d(sink0_data[86]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[5]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[5] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[5]~1 (
	.dataa(!sink0_data[68]),
	.datab(!out_data_5),
	.datac(!use_reg),
	.datad(!address_reg_5),
	.datae(!src_payload5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[5]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[5]~1 .lut_mask = 64'h101FF0FF101FF0FF;
defparam \d0_int_nxt_addr[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[5]~5 (
	.dataa(!new_burst_reg1),
	.datab(!sink0_data[86]),
	.datac(!\in_burstwrap_reg[5]~q ),
	.datad(!\int_nxt_addr_with_offset[5]~combout ),
	.datae(!\d0_int_nxt_addr[5]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[5]~5 .extended_lut = "off";
defparam \nxt_addr[5]~5 .lut_mask = 64'h00A044E400A044E4;
defparam \nxt_addr[5]~5 .shared_arith = "off";

dffeas \int_nxt_addr_reg[5] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[5]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[5]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[5] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[5] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[5] (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~21_sumout ),
	.datac(!src_data_194),
	.datad(!src_data_1941),
	.datae(!\in_burstwrap_reg[5]~q ),
	.dataf(!\int_nxt_addr_reg[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[5] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[5] .lut_mask = 64'h01112333FFFFFFFF;
defparam \int_nxt_addr_with_offset[5] .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \in_burstwrap_reg[6] (
	.clk(outclk_wire_0),
	.d(sink0_data[87]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[6]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[6] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[6]~2 (
	.dataa(!sink0_data[68]),
	.datab(!out_data_6),
	.datac(!use_reg),
	.datad(!address_reg_6),
	.datae(!src_payload6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[6]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[6]~2 .lut_mask = 64'h101FF0FF101FF0FF;
defparam \d0_int_nxt_addr[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[6]~6 (
	.dataa(!new_burst_reg1),
	.datab(!sink0_data[87]),
	.datac(!\in_burstwrap_reg[6]~q ),
	.datad(!\int_nxt_addr_with_offset[6]~combout ),
	.datae(!\d0_int_nxt_addr[6]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[6]~6 .extended_lut = "off";
defparam \nxt_addr[6]~6 .lut_mask = 64'h00A044E400A044E4;
defparam \nxt_addr[6]~6 .shared_arith = "off";

dffeas \int_nxt_addr_reg[6] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[6]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[6]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[6] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[6] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[6] (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~25_sumout ),
	.datac(!src_data_195),
	.datad(!src_data_1951),
	.datae(!\in_burstwrap_reg[6]~q ),
	.dataf(!\int_nxt_addr_reg[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[6] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[6] .lut_mask = 64'h01112333FFFFFFFF;
defparam \int_nxt_addr_with_offset[6] .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \in_burstwrap_reg[7] (
	.clk(outclk_wire_0),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[7]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[7] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[7] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[7]~3 (
	.dataa(!sink0_data[68]),
	.datab(!out_data_7),
	.datac(!use_reg),
	.datad(!address_reg_7),
	.datae(!src_payload7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[7]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[7]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[7]~3 .lut_mask = 64'h101FF0FF101FF0FF;
defparam \d0_int_nxt_addr[7]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[7]~7 (
	.dataa(!new_burst_reg1),
	.datab(!sink0_data[88]),
	.datac(!\in_burstwrap_reg[7]~q ),
	.datad(!\int_nxt_addr_with_offset[7]~combout ),
	.datae(!\d0_int_nxt_addr[7]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[7]~7 .extended_lut = "off";
defparam \nxt_addr[7]~7 .lut_mask = 64'h00A044E400A044E4;
defparam \nxt_addr[7]~7 .shared_arith = "off";

dffeas \int_nxt_addr_reg[7] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[7]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[7]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[7] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[7] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[7] (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~29_sumout ),
	.datac(!src_data_196),
	.datad(!src_data_1961),
	.datae(!\in_burstwrap_reg[7]~q ),
	.dataf(!\int_nxt_addr_reg[7]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[7] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[7] .lut_mask = 64'h01112333FFFFFFFF;
defparam \int_nxt_addr_with_offset[7] .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \in_burstwrap_reg[8] (
	.clk(outclk_wire_0),
	.d(sink0_data[89]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[8]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[8] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[8] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[8]~8 (
	.dataa(!new_burst_reg1),
	.datab(!sink0_data[89]),
	.datac(!\in_burstwrap_reg[8]~q ),
	.datad(!\int_nxt_addr_with_offset[8]~combout ),
	.datae(!out_data_44),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[8]~8 .extended_lut = "off";
defparam \nxt_addr[8]~8 .lut_mask = 64'h00A044E400A044E4;
defparam \nxt_addr[8]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg[8] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[8]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[8]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[8] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[8] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[8] (
	.dataa(!new_burst_reg1),
	.datab(!\Add0~33_sumout ),
	.datac(!src_data_197),
	.datad(!src_data_1971),
	.datae(!\in_burstwrap_reg[8]~q ),
	.dataf(!\int_nxt_addr_reg[8]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[8] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[8] .lut_mask = 64'h01112333FFFFFFFF;
defparam \int_nxt_addr_with_offset[8] .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \nxt_addr[9]~9 (
	.dataa(!new_burst_reg1),
	.datab(!sink0_data[89]),
	.datac(!\in_burstwrap_reg[8]~q ),
	.datad(!\int_nxt_addr_with_offset[9]~combout ),
	.datae(!out_data_45),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[9]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[9]~9 .extended_lut = "off";
defparam \nxt_addr[9]~9 .lut_mask = 64'h00A044E400A044E4;
defparam \nxt_addr[9]~9 .shared_arith = "off";

dffeas \int_nxt_addr_reg[9] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[9]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[9]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[9] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[9] .power_up = "low";

cyclonev_lcell_comb \int_nxt_addr_with_offset[9] (
	.dataa(!new_burst_reg1),
	.datab(!src_data_197),
	.datac(!src_data_1971),
	.datad(!\in_burstwrap_reg[8]~q ),
	.datae(!\Add0~37_sumout ),
	.dataf(!\int_nxt_addr_reg[9]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_nxt_addr_with_offset[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_nxt_addr_with_offset[9] .extended_lut = "off";
defparam \int_nxt_addr_with_offset[9] .lut_mask = 64'h000015BFFFFFFFFF;
defparam \int_nxt_addr_with_offset[9] .shared_arith = "off";

cyclonev_lcell_comb \Add4~5 (
	.dataa(!cp_ready1),
	.datab(!out_valid_reg1),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!mem_used_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~5_sumout ),
	.cout(\Add4~6 ),
	.shareout(\Add4~7 ));
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h0000EFFF00001E0F;
defparam \Add4~5 .shared_arith = "on";

cyclonev_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(\Add4~7 ),
	.combout(),
	.sumout(\Add4~9_sumout ),
	.cout(\Add4~10 ),
	.shareout(\Add4~11 ));
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h00000F0F0000F0F0;
defparam \Add4~9 .shared_arith = "on";

cyclonev_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!out_uncomp_byte_cnt_reg_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(\Add4~11 ),
	.combout(),
	.sumout(\Add4~13_sumout ),
	.cout(\Add4~14 ),
	.shareout(\Add4~15 ));
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add4~13 .shared_arith = "on";

cyclonev_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(\Add4~15 ),
	.combout(),
	.sumout(\Add4~17_sumout ),
	.cout(\Add4~18 ),
	.shareout(\Add4~19 ));
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add4~17 .shared_arith = "on";

cyclonev_lcell_comb \Add4~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!out_uncomp_byte_cnt_reg_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~18 ),
	.sharein(\Add4~19 ),
	.combout(),
	.sumout(\Add4~21_sumout ),
	.cout(\Add4~22 ),
	.shareout(\Add4~23 ));
defparam \Add4~21 .extended_lut = "off";
defparam \Add4~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add4~21 .shared_arith = "on";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~0 .lut_mask = 64'h10FE10FE10FE10FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~1 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~1 .lut_mask = 64'h10FE10FE10FE10FE;
defparam \nxt_uncomp_subburst_byte_cnt[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~2 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .lut_mask = 64'h10FE10FE10FE10FE;
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[7]~3 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[7]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[7]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[7]~3 .lut_mask = 64'h10FE10FE10FE10FE;
defparam \nxt_uncomp_subburst_byte_cnt[7]~3 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_4),
	.datae(!out_uncomp_byte_cnt_reg_8),
	.dataf(!out_uncomp_byte_cnt_reg_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hEF01010101010101;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~1 (
	.dataa(!\nxt_uncomp_subburst_byte_cnt[6]~0_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[2]~1_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[7]~3_combout ),
	.datae(!\WideOr0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~1 .extended_lut = "off";
defparam \WideOr0~1 .lut_mask = 64'h0000800000008000;
defparam \WideOr0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add4~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!out_uncomp_byte_cnt_reg_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~22 ),
	.sharein(\Add4~23 ),
	.combout(),
	.sumout(\Add4~25_sumout ),
	.cout(\Add4~26 ),
	.shareout(\Add4~27 ));
defparam \Add4~25 .extended_lut = "off";
defparam \Add4~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add4~25 .shared_arith = "on";

cyclonev_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!out_uncomp_byte_cnt_reg_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~26 ),
	.sharein(\Add4~27 ),
	.combout(),
	.sumout(\Add4~1_sumout ),
	.cout(),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h000000000000FF00;
defparam \Add4~1 .shared_arith = "on";

cyclonev_lcell_comb \WideOr0~2 (
	.dataa(!\Add4~5_sumout ),
	.datab(!\Add4~9_sumout ),
	.datac(!\Add4~13_sumout ),
	.datad(!\Add4~17_sumout ),
	.datae(!\Add4~21_sumout ),
	.dataf(!\Add4~25_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~2 .extended_lut = "off";
defparam \WideOr0~2 .lut_mask = 64'h8000000000000000;
defparam \WideOr0~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_in_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h8888888888888888;
defparam \nxt_in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!cp_ready),
	.datac(!in_eop_reg1),
	.datad(!new_burst_reg1),
	.datae(!in_bytecount_reg_zero1),
	.dataf(!\nxt_in_ready~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'hF5E4B1A000000000;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!in_ready_hold),
	.datab(!source0_data_33),
	.datac(!WideOr0),
	.datad(!mem_used_1),
	.datae(!new_burst_reg1),
	.dataf(!in_bytecount_reg_zero1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_eop~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h00005D00A2FFFFFF;
defparam \nxt_out_eop~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[69]),
	.datac(!sink0_data[68]),
	.datad(!nxt_out_eop),
	.datae(!WideOr1),
	.dataf(!\state.ST_IDLE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h00001515FF00FF55;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(outclk_wire_0),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_eop_reg1),
	.datac(!\nxt_out_eop~0_combout ),
	.datad(!stateST_UNCOMP_WR_SUBBURST),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h0000FAD80000FAD8;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!in_ready_hold),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!WideOr1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0101010101010101;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[69]),
	.datac(!nxt_out_eop),
	.datad(!src_valid),
	.datae(!\Selector2~0_combout ),
	.dataf(!\Selector2~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "off";
defparam \Selector2~2 .lut_mask = 64'h004400000C4C0C0C;
defparam \Selector2~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\WideOr0~1_combout ),
	.datac(!\Add4~1_sumout ),
	.datad(!\WideOr0~2_combout ),
	.datae(!\Selector3~0_combout ),
	.dataf(!\Selector2~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~3 .extended_lut = "off";
defparam \Selector2~3 .lut_mask = 64'h000011B1FFFFFFFF;
defparam \Selector2~3 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(outclk_wire_0),
	.d(\Selector2~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~4 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .lut_mask = 64'h10FE10FE10FE10FE;
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[8]~5 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[8]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[8]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[8]~5 .lut_mask = 64'h10FE10FE10FE10FE;
defparam \nxt_uncomp_subburst_byte_cnt[8]~5 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~6 (
	.dataa(!out_valid_reg1),
	.datab(!cp_ready),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~6 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~6 .lut_mask = 64'h10FE10FE10FE10FE;
defparam \nxt_uncomp_subburst_byte_cnt[5]~6 .shared_arith = "off";

cyclonev_lcell_comb \always10~0 (
	.dataa(!out_valid_reg1),
	.datab(!stateST_COMP_TRANS),
	.datac(!cp_ready),
	.datad(gnd),
	.datae(!new_burst_reg1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~0 .extended_lut = "off";
defparam \always10~0 .lut_mask = 64'hAEAEAFAFAEAEAFAF;
defparam \always10~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!sink0_data[69]),
	.datab(!stateST_COMP_TRANS),
	.datac(!in_eop_reg1),
	.datad(!\nxt_in_ready~1_combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h5555151155551511;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[68]),
	.datac(!stateST_COMP_TRANS),
	.datad(!nxt_out_eop),
	.datae(!WideOr1),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h0F000F040F005F55;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \in_narrow_reg~0 (
	.dataa(!sink0_data[91]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_narrow_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_narrow_reg~0 .extended_lut = "off";
defparam \in_narrow_reg~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \in_narrow_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!out_data_79),
	.datab(!out_data_76),
	.datac(!out_data_77),
	.datad(!out_data_78),
	.datae(!out_data_80),
	.dataf(!out_data_75),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'h8000000000000000;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(outclk_wire_0),
	.d(\Add1~1_sumout ),
	.asdata(out_data_77),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout(\Add1~19 ));
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add1~17 .shared_arith = "on";

dffeas \int_bytes_remaining_reg[2] (
	.clk(outclk_wire_0),
	.d(\Add1~17_sumout ),
	.asdata(out_data_74),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(\Add1~19 ),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout(\Add1~23 ));
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add1~21 .shared_arith = "on";

dffeas \int_bytes_remaining_reg[3] (
	.clk(outclk_wire_0),
	.d(\Add1~21_sumout ),
	.asdata(out_data_75),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_bytes_remaining_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(\Add1~23 ),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout(\Add1~27 ));
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add1~25 .shared_arith = "on";

dffeas \int_bytes_remaining_reg[4] (
	.clk(outclk_wire_0),
	.d(\Add1~25_sumout ),
	.asdata(out_data_76),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(\Add1~27 ),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout(\Add1~3 ));
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h000000FF0000FF00;
defparam \Add1~1 .shared_arith = "on";

dffeas \int_bytes_remaining_reg[6] (
	.clk(outclk_wire_0),
	.d(\Add1~5_sumout ),
	.asdata(out_data_78),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_bytes_remaining_reg[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(\Add1~3 ),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout(\Add1~7 ));
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add1~5 .shared_arith = "on";

dffeas \int_bytes_remaining_reg[7] (
	.clk(outclk_wire_0),
	.d(\Add1~9_sumout ),
	.asdata(out_data_79),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[7]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[7] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[7] .power_up = "low";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_bytes_remaining_reg[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(\Add1~7 ),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout(\Add1~11 ));
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add1~9 .shared_arith = "on";

dffeas \int_bytes_remaining_reg[8] (
	.clk(outclk_wire_0),
	.d(\Add1~13_sumout ),
	.asdata(out_data_80),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(new_burst_reg1),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[8]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[8] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[8] .power_up = "low";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_bytes_remaining_reg[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(\Add1~11 ),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h000000000000FF00;
defparam \Add1~13 .shared_arith = "on";

cyclonev_lcell_comb \new_burst_reg~1 (
	.dataa(!new_burst_reg1),
	.datab(!\Add1~17_sumout ),
	.datac(!\Add1~21_sumout ),
	.datad(!\Add1~25_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~1 .extended_lut = "off";
defparam \new_burst_reg~1 .lut_mask = 64'h2000200020002000;
defparam \new_burst_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~2 (
	.dataa(!\Add1~1_sumout ),
	.datab(!\Add1~5_sumout ),
	.datac(!\Add1~9_sumout ),
	.datad(!\Add1~13_sumout ),
	.datae(!\new_burst_reg~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~2 .extended_lut = "off";
defparam \new_burst_reg~2 .lut_mask = 64'h0000800000008000;
defparam \new_burst_reg~2 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~3 (
	.dataa(!new_burst_reg1),
	.datab(!\Selector1~1_combout ),
	.datac(!out_data_74),
	.datad(!\new_burst_reg~0_combout ),
	.datae(!\new_burst_reg~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~3 .extended_lut = "off";
defparam \new_burst_reg~3 .lut_mask = 64'hCCCDFFFFCCCDFFFF;
defparam \new_burst_reg~3 .shared_arith = "off";

cyclonev_lcell_comb WideNor0(
	.dataa(!out_data_74),
	.datab(!\new_burst_reg~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor0.extended_lut = "off";
defparam WideNor0.lut_mask = 64'h2222222222222222;
defparam WideNor0.shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!in_bytecount_reg_zero1),
	.datab(!new_burst_reg1),
	.datac(!WideOr1),
	.datad(!mem_used_1),
	.datae(!in_ready_hold),
	.dataf(!stateST_COMP_TRANS),
	.datag(!cp_ready2),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "on";
defparam \nxt_out_valid~0 .lut_mask = 64'h00000F0FACAACFAF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~3 (
	.dataa(!\Add4~5_sumout ),
	.datab(!\Add4~9_sumout ),
	.datac(!\Add4~13_sumout ),
	.datad(!\Add4~17_sumout ),
	.datae(!\Add4~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~3 .extended_lut = "off";
defparam \WideOr0~3 .lut_mask = 64'h8000000080000000;
defparam \WideOr0~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\WideOr0~1_combout ),
	.datac(!\Add4~25_sumout ),
	.datad(!\Add4~1_sumout ),
	.datae(!\WideOr0~3_combout ),
	.dataf(!\Selector3~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~1 .extended_lut = "off";
defparam \Selector3~1 .lut_mask = 64'h00000000EEEE4EEE;
defparam \Selector3~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~3 (
	.dataa(!in_ready_hold),
	.datab(!out_valid_reg1),
	.datac(!source0_data_33),
	.datad(!WideOr0),
	.datae(!mem_used_1),
	.dataf(!\nxt_in_ready~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_in_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~3 .extended_lut = "off";
defparam \nxt_in_ready~3 .lut_mask = 64'h22023333AAAAAAAA;
defparam \nxt_in_ready~3 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_address_alignment_2 (
	src_data_198,
	src_data_199,
	src_data_200,
	in_data_reg_91,
	in_data_reg_90,
	new_burst_reg,
	out_data_91,
	out_data_37,
	out_data_1,
	LessThan0,
	out_data_36,
	out_data_0)/* synthesis synthesis_greybox=0 */;
input 	src_data_198;
input 	src_data_199;
input 	src_data_200;
input 	in_data_reg_91;
input 	in_data_reg_90;
input 	new_burst_reg;
input 	out_data_91;
input 	out_data_37;
output 	out_data_1;
output 	LessThan0;
input 	out_data_36;
output 	out_data_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \out_data[1] (
	.dataa(!in_data_reg_91),
	.datab(!new_burst_reg),
	.datac(!out_data_91),
	.datad(!out_data_37),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[1] .extended_lut = "off";
defparam \out_data[1] .lut_mask = 64'h00B800B800B800B8;
defparam \out_data[1] .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!src_data_198),
	.datab(!src_data_199),
	.datac(!src_data_200),
	.datad(!in_data_reg_91),
	.datae(!in_data_reg_90),
	.dataf(!new_burst_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hFF00000080808080;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[0] (
	.dataa(!LessThan0),
	.datab(!out_data_36),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[0] .extended_lut = "off";
defparam \out_data[0] .lut_mask = 64'h1111111111111111;
defparam \out_data[0] .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_slave_agent (
	outclk_wire_0,
	op_2,
	op_21,
	op_22,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wrfull,
	wrfull1,
	mem_used_1,
	mem_125_0,
	mem_used_0,
	comb,
	mem_90_0,
	mem_91_0,
	mem_38_0,
	source_addr_2,
	mem_39_0,
	source_addr_3,
	in_data_reg_68,
	nxt_uncomp_subburst_byte_cnt,
	m0_write,
	r_sync_rst,
	wrfull2,
	cp_ready,
	read,
	cp_ready1,
	mem_83_0,
	mem_84_0,
	mem_37_0,
	mem_82_0,
	mem_36_0,
	mem_81_0)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
input 	op_2;
input 	op_21;
input 	op_22;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wrfull;
input 	wrfull1;
input 	mem_used_1;
input 	mem_125_0;
input 	mem_used_0;
output 	comb;
input 	mem_90_0;
input 	mem_91_0;
input 	mem_38_0;
output 	source_addr_2;
input 	mem_39_0;
output 	source_addr_3;
input 	in_data_reg_68;
input 	nxt_uncomp_subburst_byte_cnt;
output 	m0_write;
input 	r_sync_rst;
input 	wrfull2;
output 	cp_ready;
input 	read;
output 	cp_ready1;
input 	mem_83_0;
input 	mem_84_0;
input 	mem_37_0;
input 	mem_82_0;
input 	mem_36_0;
input 	mem_81_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altera_merlin_burst_uncompressor uncompressor(
	.clk(outclk_wire_0),
	.mem_125_0(mem_125_0),
	.mem_used_0(mem_used_0),
	.mem_90_0(mem_90_0),
	.mem_91_0(mem_91_0),
	.mem_38_0(mem_38_0),
	.source_addr_2(source_addr_2),
	.mem_39_0(mem_39_0),
	.source_addr_3(source_addr_3),
	.reset(r_sync_rst),
	.read(read),
	.mem_83_0(mem_83_0),
	.mem_84_0(mem_84_0),
	.mem_37_0(mem_37_0),
	.mem_82_0(mem_82_0),
	.mem_36_0(mem_36_0),
	.mem_81_0(mem_81_0));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h8000800080008000;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!mem_125_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h1111111111111111;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb \m0_write~0 (
	.dataa(!WideOr0),
	.datab(!in_data_reg_68),
	.datac(!nxt_uncomp_subburst_byte_cnt),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'h0202020202020202;
defparam \m0_write~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!op_2),
	.datab(!op_21),
	.datac(!op_22),
	.datad(!WideOr0),
	.datae(!wrfull2),
	.dataf(!wrfull1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'h00FF00FFFFFFFEFF;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!op_21),
	.datab(!op_22),
	.datac(!WideOr0),
	.datad(!wrfull),
	.datae(!wrfull1),
	.dataf(!mem_used_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h0F0FFFEF00000000;
defparam \cp_ready~1 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_burst_uncompressor (
	clk,
	mem_125_0,
	mem_used_0,
	mem_90_0,
	mem_91_0,
	mem_38_0,
	source_addr_2,
	mem_39_0,
	source_addr_3,
	reset,
	read,
	mem_83_0,
	mem_84_0,
	mem_37_0,
	mem_82_0,
	mem_36_0,
	mem_81_0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	mem_125_0;
input 	mem_used_0;
input 	mem_90_0;
input 	mem_91_0;
input 	mem_38_0;
output 	source_addr_2;
input 	mem_39_0;
output 	source_addr_3;
input 	reset;
input 	read;
input 	mem_83_0;
input 	mem_84_0;
input 	mem_37_0;
input 	mem_82_0;
input 	mem_36_0;
input 	mem_81_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_address_base~0_combout ;
wire \burst_uncompress_address_base[2]~q ;
wire \Decoder0~0_combout ;
wire \Decoder0~2_combout ;
wire \Decoder0~3_combout ;
wire \Add2~13_sumout ;
wire \p1_burst_uncompress_address_offset[0]~combout ;
wire \burst_uncompress_address_offset[0]~q ;
wire \Add2~14 ;
wire \Add2~9_sumout ;
wire \p1_burst_uncompress_address_offset[1]~combout ;
wire \burst_uncompress_address_offset[1]~q ;
wire \Add2~10 ;
wire \Add2~1_sumout ;
wire \p1_burst_uncompress_address_offset[2]~combout ;
wire \burst_uncompress_address_offset[2]~q ;
wire \burst_uncompress_address_base~1_combout ;
wire \burst_uncompress_address_base[3]~q ;
wire \Decoder0~1_combout ;
wire \Add2~2 ;
wire \Add2~5_sumout ;
wire \p1_burst_uncompress_address_offset[3]~combout ;
wire \burst_uncompress_address_offset[3]~q ;


cyclonev_lcell_comb \source_addr[2]~0 (
	.dataa(!mem_38_0),
	.datab(!mem_125_0),
	.datac(!mem_used_0),
	.datad(!\burst_uncompress_address_base[2]~q ),
	.datae(!\burst_uncompress_address_offset[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_addr_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_addr[2]~0 .extended_lut = "off";
defparam \source_addr[2]~0 .lut_mask = 64'hFE020202FE020202;
defparam \source_addr[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \source_addr[3]~1 (
	.dataa(!mem_125_0),
	.datab(!mem_used_0),
	.datac(!mem_39_0),
	.datad(!\burst_uncompress_address_base[3]~q ),
	.datae(!\burst_uncompress_address_offset[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_addr_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_addr[3]~1 .extended_lut = "off";
defparam \source_addr[3]~1 .lut_mask = 64'hFE101010FE101010;
defparam \source_addr[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_address_base~0 (
	.dataa(!mem_38_0),
	.datab(!mem_83_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_address_base~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_address_base~0 .extended_lut = "off";
defparam \burst_uncompress_address_base~0 .lut_mask = 64'h4444444444444444;
defparam \burst_uncompress_address_base~0 .shared_arith = "off";

dffeas \burst_uncompress_address_base[2] (
	.clk(clk),
	.d(\burst_uncompress_address_base~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_address_base[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_base[2] .is_wysiwyg = "true";
defparam \burst_uncompress_address_base[2] .power_up = "low";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!mem_90_0),
	.datab(!mem_91_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'h2222222222222222;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~2 (
	.dataa(!mem_90_0),
	.datab(!mem_91_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~2 .extended_lut = "off";
defparam \Decoder0~2 .lut_mask = 64'h4444444444444444;
defparam \Decoder0~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~3 (
	.dataa(!mem_90_0),
	.datab(!mem_91_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~3 .extended_lut = "off";
defparam \Decoder0~3 .lut_mask = 64'h8888888888888888;
defparam \Decoder0~3 .shared_arith = "off";

cyclonev_lcell_comb \Add2~13 (
	.dataa(!mem_125_0),
	.datab(!mem_used_0),
	.datac(!mem_36_0),
	.datad(!\Decoder0~3_combout ),
	.datae(gnd),
	.dataf(!\burst_uncompress_address_offset[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h0000FE10000000FF;
defparam \Add2~13 .shared_arith = "off";

cyclonev_lcell_comb \p1_burst_uncompress_address_offset[0] (
	.dataa(!\Add2~13_sumout ),
	.datab(!mem_81_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_burst_uncompress_address_offset[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_burst_uncompress_address_offset[0] .extended_lut = "off";
defparam \p1_burst_uncompress_address_offset[0] .lut_mask = 64'h1111111111111111;
defparam \p1_burst_uncompress_address_offset[0] .shared_arith = "off";

dffeas \burst_uncompress_address_offset[0] (
	.clk(clk),
	.d(\p1_burst_uncompress_address_offset[0]~combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_address_offset[0]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_offset[0] .is_wysiwyg = "true";
defparam \burst_uncompress_address_offset[0] .power_up = "low";

cyclonev_lcell_comb \Add2~9 (
	.dataa(!mem_125_0),
	.datab(!mem_used_0),
	.datac(!mem_37_0),
	.datad(!\Decoder0~2_combout ),
	.datae(gnd),
	.dataf(!\burst_uncompress_address_offset[1]~q ),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h0000FE10000000FF;
defparam \Add2~9 .shared_arith = "off";

cyclonev_lcell_comb \p1_burst_uncompress_address_offset[1] (
	.dataa(!\Add2~9_sumout ),
	.datab(!mem_82_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_burst_uncompress_address_offset[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_burst_uncompress_address_offset[1] .extended_lut = "off";
defparam \p1_burst_uncompress_address_offset[1] .lut_mask = 64'h1111111111111111;
defparam \p1_burst_uncompress_address_offset[1] .shared_arith = "off";

dffeas \burst_uncompress_address_offset[1] (
	.clk(clk),
	.d(\p1_burst_uncompress_address_offset[1]~combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_address_offset[1]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_offset[1] .is_wysiwyg = "true";
defparam \burst_uncompress_address_offset[1] .power_up = "low";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!mem_125_0),
	.datab(!mem_used_0),
	.datac(!mem_38_0),
	.datad(!\Decoder0~0_combout ),
	.datae(gnd),
	.dataf(!\burst_uncompress_address_offset[2]~q ),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h0000FE10000000FF;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_burst_uncompress_address_offset[2] (
	.dataa(!mem_83_0),
	.datab(!\Add2~1_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_burst_uncompress_address_offset[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_burst_uncompress_address_offset[2] .extended_lut = "off";
defparam \p1_burst_uncompress_address_offset[2] .lut_mask = 64'h1111111111111111;
defparam \p1_burst_uncompress_address_offset[2] .shared_arith = "off";

dffeas \burst_uncompress_address_offset[2] (
	.clk(clk),
	.d(\p1_burst_uncompress_address_offset[2]~combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_address_offset[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_offset[2] .is_wysiwyg = "true";
defparam \burst_uncompress_address_offset[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_address_base~1 (
	.dataa(!mem_39_0),
	.datab(!mem_84_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_address_base~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_address_base~1 .extended_lut = "off";
defparam \burst_uncompress_address_base~1 .lut_mask = 64'h4444444444444444;
defparam \burst_uncompress_address_base~1 .shared_arith = "off";

dffeas \burst_uncompress_address_base[3] (
	.clk(clk),
	.d(\burst_uncompress_address_base~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_address_base[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_base[3] .is_wysiwyg = "true";
defparam \burst_uncompress_address_base[3] .power_up = "low";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!mem_90_0),
	.datab(!mem_91_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'h1111111111111111;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add2~5 (
	.dataa(!mem_125_0),
	.datab(!mem_used_0),
	.datac(!mem_39_0),
	.datad(!\Decoder0~1_combout ),
	.datae(gnd),
	.dataf(!\burst_uncompress_address_offset[3]~q ),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h0000FE10000000FF;
defparam \Add2~5 .shared_arith = "off";

cyclonev_lcell_comb \p1_burst_uncompress_address_offset[3] (
	.dataa(!mem_84_0),
	.datab(!\Add2~5_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_burst_uncompress_address_offset[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_burst_uncompress_address_offset[3] .extended_lut = "off";
defparam \p1_burst_uncompress_address_offset[3] .lut_mask = 64'h1111111111111111;
defparam \p1_burst_uncompress_address_offset[3] .shared_arith = "off";

dffeas \burst_uncompress_address_offset[3] (
	.clk(clk),
	.d(\p1_burst_uncompress_address_offset[3]~combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_address_offset[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_offset[3] .is_wysiwyg = "true";
defparam \burst_uncompress_address_offset[3] .power_up = "low";

endmodule

module Computer_System_altera_merlin_slave_agent_1 (
	outclk_wire_0,
	in_ready_hold,
	in_narrow_reg,
	always12,
	in_byteen_reg_2,
	source0_data_34,
	in_byteen_reg_0,
	source0_data_32,
	in_byteen_reg_1,
	source0_data_33,
	in_byteen_reg_3,
	source0_data_35,
	source0_data_351,
	mem_used_1,
	cp_ready1,
	out_valid_reg,
	ShiftLeft1,
	source0_data_352,
	WideOr01,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_125_0,
	mem_used_01,
	out_valid,
	comb,
	mem_66_0,
	burst_uncompress_busy,
	last_packet_beat,
	last_packet_beat1,
	mem_80_0,
	mem_79_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat2,
	src_payload,
	mem_38_0,
	source_addr_2,
	source_addr_21,
	mem_91_0,
	mem_90_0,
	mem_39_0,
	source_addr_3,
	always10,
	in_data_reg_68,
	m0_write,
	r_sync_rst,
	last_packet_beat3,
	p1_ready,
	cp_ready2,
	cp_ready3,
	WideOr02,
	mem_83_0,
	mem_84_0,
	mem_37_0,
	mem_82_0,
	mem_36_0,
	mem_81_0)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
input 	in_ready_hold;
input 	in_narrow_reg;
input 	always12;
input 	in_byteen_reg_2;
input 	source0_data_34;
input 	in_byteen_reg_0;
input 	source0_data_32;
input 	in_byteen_reg_1;
input 	source0_data_33;
input 	in_byteen_reg_3;
input 	source0_data_35;
input 	source0_data_351;
input 	mem_used_1;
output 	cp_ready1;
input 	out_valid_reg;
input 	ShiftLeft1;
input 	source0_data_352;
output 	WideOr01;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_125_0;
input 	mem_used_01;
input 	out_valid;
output 	comb;
input 	mem_66_0;
output 	burst_uncompress_busy;
output 	last_packet_beat;
output 	last_packet_beat1;
input 	mem_80_0;
input 	mem_79_0;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat2;
input 	src_payload;
input 	mem_38_0;
output 	source_addr_2;
output 	source_addr_21;
input 	mem_91_0;
input 	mem_90_0;
input 	mem_39_0;
output 	source_addr_3;
input 	always10;
input 	in_data_reg_68;
output 	m0_write;
input 	r_sync_rst;
output 	last_packet_beat3;
input 	p1_ready;
output 	cp_ready2;
output 	cp_ready3;
output 	WideOr02;
input 	mem_83_0;
input 	mem_84_0;
input 	mem_37_0;
input 	mem_82_0;
input 	mem_36_0;
input 	mem_81_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altera_merlin_burst_uncompressor_1 uncompressor(
	.clk(outclk_wire_0),
	.out_valid(out_valid),
	.comb(comb),
	.mem_66_0(mem_66_0),
	.burst_uncompress_busy1(burst_uncompress_busy),
	.last_packet_beat(last_packet_beat),
	.last_packet_beat1(last_packet_beat1),
	.mem_80_0(mem_80_0),
	.mem_79_0(mem_79_0),
	.mem_78_0(mem_78_0),
	.mem_77_0(mem_77_0),
	.mem_76_0(mem_76_0),
	.mem_75_0(mem_75_0),
	.mem_74_0(mem_74_0),
	.last_packet_beat2(last_packet_beat2),
	.src_payload(src_payload),
	.mem_38_0(mem_38_0),
	.source_addr_2(source_addr_2),
	.source_addr_21(source_addr_21),
	.mem_91_0(mem_91_0),
	.mem_90_0(mem_90_0),
	.mem_39_0(mem_39_0),
	.source_addr_3(source_addr_3),
	.always10(always10),
	.reset(r_sync_rst),
	.last_packet_beat3(last_packet_beat3),
	.p1_ready(p1_ready),
	.mem_83_0(mem_83_0),
	.mem_84_0(mem_84_0),
	.mem_37_0(mem_37_0),
	.mem_82_0(mem_82_0),
	.mem_36_0(mem_36_0),
	.mem_81_0(mem_81_0));

cyclonev_lcell_comb cp_ready(
	.dataa(!in_ready_hold),
	.datab(!source0_data_34),
	.datac(!source0_data_32),
	.datad(!source0_data_33),
	.datae(!source0_data_351),
	.dataf(!mem_used_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam cp_ready.extended_lut = "off";
defparam cp_ready.lut_mask = 64'hD555555500000000;
defparam cp_ready.shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!always12),
	.datab(!ShiftLeft1),
	.datac(!in_byteen_reg_2),
	.datad(!source0_data_32),
	.datae(!source0_data_352),
	.dataf(!source0_data_35),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr01),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hB100000000000000;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_125_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb \m0_write~0 (
	.dataa(!out_valid_reg),
	.datab(!source0_data_33),
	.datac(!WideOr01),
	.datad(!mem_used_1),
	.datae(!in_data_reg_68),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'h0000510000005100;
defparam \m0_write~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!in_ready_hold),
	.datab(!source0_data_34),
	.datac(!source0_data_32),
	.datad(!source0_data_33),
	.datae(!source0_data_351),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hD5555555D5555555;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_narrow_reg),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_0),
	.datad(!in_byteen_reg_1),
	.datae(!in_byteen_reg_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready3),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000000080000000;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!source0_data_34),
	.datab(!source0_data_32),
	.datac(!source0_data_33),
	.datad(!source0_data_351),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr02),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h8000800080008000;
defparam WideOr0.shared_arith = "off";

endmodule

module Computer_System_altera_merlin_burst_uncompressor_1 (
	clk,
	out_valid,
	comb,
	mem_66_0,
	burst_uncompress_busy1,
	last_packet_beat,
	last_packet_beat1,
	mem_80_0,
	mem_79_0,
	mem_78_0,
	mem_77_0,
	mem_76_0,
	mem_75_0,
	mem_74_0,
	last_packet_beat2,
	src_payload,
	mem_38_0,
	source_addr_2,
	source_addr_21,
	mem_91_0,
	mem_90_0,
	mem_39_0,
	source_addr_3,
	always10,
	reset,
	last_packet_beat3,
	p1_ready,
	mem_83_0,
	mem_84_0,
	mem_37_0,
	mem_82_0,
	mem_36_0,
	mem_81_0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	out_valid;
input 	comb;
input 	mem_66_0;
output 	burst_uncompress_busy1;
output 	last_packet_beat;
output 	last_packet_beat1;
input 	mem_80_0;
input 	mem_79_0;
input 	mem_78_0;
input 	mem_77_0;
input 	mem_76_0;
input 	mem_75_0;
input 	mem_74_0;
output 	last_packet_beat2;
input 	src_payload;
input 	mem_38_0;
output 	source_addr_2;
output 	source_addr_21;
input 	mem_91_0;
input 	mem_90_0;
input 	mem_39_0;
output 	source_addr_3;
input 	always10;
input 	reset;
output 	last_packet_beat3;
input 	p1_ready;
input 	mem_83_0;
input 	mem_84_0;
input 	mem_37_0;
input 	mem_82_0;
input 	mem_36_0;
input 	mem_81_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~0_combout ;
wire \burst_uncompress_busy~0_combout ;
wire \Add0~30_cout ;
wire \Add0~17_sumout ;
wire \Add1~30_cout ;
wire \Add1~17_sumout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \burst_uncompress_byte_counter~7_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \Add0~22 ;
wire \Add0~13_sumout ;
wire \Add1~22 ;
wire \Add1~13_sumout ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \Add1~14 ;
wire \Add1~9_sumout ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[6]~q ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \Add1~10 ;
wire \Add1~5_sumout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \Add1~6 ;
wire \Add1~1_sumout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[8]~q ;
wire \Add0~2 ;
wire \Add0~25_sumout ;
wire \Add1~2 ;
wire \Add1~25_sumout ;
wire \burst_uncompress_byte_counter~8_combout ;
wire \burst_uncompress_byte_counter[9]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \last_packet_beat~2_combout ;
wire \last_packet_beat~3_combout ;
wire \burst_uncompress_address_base~0_combout ;
wire \always1~0_combout ;
wire \burst_uncompress_address_base[2]~q ;
wire \Decoder0~0_combout ;
wire \Decoder0~2_combout ;
wire \Decoder0~3_combout ;
wire \Add2~13_sumout ;
wire \p1_burst_uncompress_address_offset[0]~combout ;
wire \burst_uncompress_address_offset[0]~q ;
wire \Add2~14 ;
wire \Add2~9_sumout ;
wire \p1_burst_uncompress_address_offset[1]~combout ;
wire \burst_uncompress_address_offset[1]~q ;
wire \Add2~10 ;
wire \Add2~1_sumout ;
wire \p1_burst_uncompress_address_offset[2]~combout ;
wire \burst_uncompress_address_offset[2]~q ;
wire \burst_uncompress_address_base~1_combout ;
wire \burst_uncompress_address_base[3]~q ;
wire \Decoder0~1_combout ;
wire \Add2~2 ;
wire \Add2~5_sumout ;
wire \p1_burst_uncompress_address_offset[3]~combout ;
wire \burst_uncompress_address_offset[3]~q ;


dffeas burst_uncompress_busy(
	.clk(clk),
	.d(\burst_uncompress_busy~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(burst_uncompress_busy1),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!burst_uncompress_busy1),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h1111111111111111;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_byte_counter[8]~q ),
	.datab(!\burst_uncompress_byte_counter[7]~q ),
	.datac(!\burst_uncompress_byte_counter[6]~q ),
	.datad(!\burst_uncompress_byte_counter[5]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h8000000000000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~4 (
	.dataa(!\last_packet_beat~2_combout ),
	.datab(!\last_packet_beat~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~4 .extended_lut = "off";
defparam \last_packet_beat~4 .lut_mask = 64'h1111111111111111;
defparam \last_packet_beat~4 .shared_arith = "off";

cyclonev_lcell_comb \source_addr[2]~0 (
	.dataa(!\burst_uncompress_address_base[2]~q ),
	.datab(!\burst_uncompress_address_offset[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_addr_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_addr[2]~0 .extended_lut = "off";
defparam \source_addr[2]~0 .lut_mask = 64'h8888888888888888;
defparam \source_addr[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \source_addr[2]~1 (
	.dataa(!comb),
	.datab(!burst_uncompress_busy1),
	.datac(!mem_38_0),
	.datad(!source_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_addr_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_addr[2]~1 .extended_lut = "off";
defparam \source_addr[2]~1 .lut_mask = 64'hBF04BF04BF04BF04;
defparam \source_addr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \source_addr[3]~2 (
	.dataa(!\burst_uncompress_address_base[3]~q ),
	.datab(!\burst_uncompress_address_offset[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_addr_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_addr[3]~2 .extended_lut = "off";
defparam \source_addr[3]~2 .lut_mask = 64'h8888888888888888;
defparam \source_addr[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~5 (
	.dataa(!comb),
	.datab(!mem_66_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(!\last_packet_beat~2_combout ),
	.dataf(!\last_packet_beat~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat3),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~5 .extended_lut = "off";
defparam \last_packet_beat~5 .lut_mask = 64'hCCCDCCCDCCCDDDDD;
defparam \last_packet_beat~5 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!comb),
	.datab(!out_valid),
	.datac(!src_payload),
	.datad(!always10),
	.datae(!p1_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h1151555511515555;
defparam \sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_busy~0 (
	.dataa(!burst_uncompress_busy1),
	.datab(!last_packet_beat3),
	.datac(!\sink_ready~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_busy~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_busy~0 .extended_lut = "off";
defparam \burst_uncompress_busy~0 .lut_mask = 64'h5C5C5C5C5C5C5C5C;
defparam \burst_uncompress_busy~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~30 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~30_cout ),
	.shareout());
defparam \Add0~30 .extended_lut = "off";
defparam \Add0~30 .lut_mask = 64'h00000000000000FF;
defparam \Add0~30 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~30 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!mem_74_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add1~30_cout ),
	.shareout());
defparam \Add1~30 .extended_lut = "off";
defparam \Add1~30 .lut_mask = 64'h00000000000000FF;
defparam \Add1~30 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!mem_75_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~30_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h00000000000000FF;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!\burst_uncompress_byte_counter~0_combout ),
	.datab(!\Add0~17_sumout ),
	.datac(!\Add1~17_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(last_packet_beat3),
	.sload(gnd),
	.ena(\sink_ready~0_combout ),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!mem_76_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h00000000000000FF;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~7 (
	.dataa(!\burst_uncompress_byte_counter~0_combout ),
	.datab(!\Add0~21_sumout ),
	.datac(!\Add1~21_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~7 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \burst_uncompress_byte_counter~7 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(last_packet_beat3),
	.sload(gnd),
	.ena(\sink_ready~0_combout ),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\burst_uncompress_byte_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!mem_77_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h00000000000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_byte_counter~0_combout ),
	.datab(!\Add0~13_sumout ),
	.datac(!\Add1~13_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(last_packet_beat3),
	.sload(gnd),
	.ena(\sink_ready~0_combout ),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\burst_uncompress_byte_counter[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!mem_78_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h00000000000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!\burst_uncompress_byte_counter~0_combout ),
	.datab(!\Add0~9_sumout ),
	.datac(!\Add1~9_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(last_packet_beat3),
	.sload(gnd),
	.ena(\sink_ready~0_combout ),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!mem_79_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h00000000000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!\burst_uncompress_byte_counter~0_combout ),
	.datab(!\Add0~5_sumout ),
	.datac(!\Add1~5_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(last_packet_beat3),
	.sload(gnd),
	.ena(\sink_ready~0_combout ),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\burst_uncompress_byte_counter[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!mem_80_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h00000000000000FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!\burst_uncompress_byte_counter~0_combout ),
	.datab(!\Add0~1_sumout ),
	.datac(!\Add1~1_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[8] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(last_packet_beat3),
	.sload(gnd),
	.ena(\sink_ready~0_combout ),
	.q(\burst_uncompress_byte_counter[8]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[8] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[8] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FFFF0000FFFF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h0000FFFF0000FFFF;
defparam \Add1~25 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~8 (
	.dataa(!\burst_uncompress_byte_counter~0_combout ),
	.datab(!\Add0~25_sumout ),
	.datac(!\Add1~25_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~8 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \burst_uncompress_byte_counter~8 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[9] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(last_packet_beat3),
	.sload(gnd),
	.ena(\sink_ready~0_combout ),
	.q(\burst_uncompress_byte_counter[9]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[9] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[9] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!burst_uncompress_busy1),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!last_packet_beat1),
	.datad(!\burst_uncompress_byte_counter[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!last_packet_beat),
	.datab(!mem_74_0),
	.datac(!\burst_uncompress_byte_counter~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(last_packet_beat3),
	.sload(gnd),
	.ena(\sink_ready~0_combout ),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!burst_uncompress_busy1),
	.datab(!mem_80_0),
	.datac(!mem_79_0),
	.datad(!mem_78_0),
	.datae(!mem_77_0),
	.dataf(!mem_76_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h8000000000000000;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!mem_75_0),
	.datab(!mem_74_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h2222222222222222;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_address_base~0 (
	.dataa(!mem_38_0),
	.datab(!mem_83_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_address_base~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_address_base~0 .extended_lut = "off";
defparam \burst_uncompress_address_base~0 .lut_mask = 64'h4444444444444444;
defparam \burst_uncompress_address_base~0 .shared_arith = "off";

cyclonev_lcell_comb \always1~0 (
	.dataa(!comb),
	.datab(!out_valid),
	.datac(!burst_uncompress_busy1),
	.datad(!src_payload),
	.datae(!always10),
	.dataf(!p1_ready),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'h1010501050505050;
defparam \always1~0 .shared_arith = "off";

dffeas \burst_uncompress_address_base[2] (
	.clk(clk),
	.d(\burst_uncompress_address_base~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\burst_uncompress_address_base[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_base[2] .is_wysiwyg = "true";
defparam \burst_uncompress_address_base[2] .power_up = "low";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!mem_90_0),
	.datab(!mem_91_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'h2222222222222222;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~2 (
	.dataa(!mem_90_0),
	.datab(!mem_91_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~2 .extended_lut = "off";
defparam \Decoder0~2 .lut_mask = 64'h4444444444444444;
defparam \Decoder0~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~3 (
	.dataa(!mem_90_0),
	.datab(!mem_91_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~3 .extended_lut = "off";
defparam \Decoder0~3 .lut_mask = 64'h8888888888888888;
defparam \Decoder0~3 .shared_arith = "off";

cyclonev_lcell_comb \Add2~13 (
	.dataa(!comb),
	.datab(!burst_uncompress_busy1),
	.datac(!mem_36_0),
	.datad(!\Decoder0~3_combout ),
	.datae(gnd),
	.dataf(!\burst_uncompress_address_offset[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h0000FB40000000FF;
defparam \Add2~13 .shared_arith = "off";

cyclonev_lcell_comb \p1_burst_uncompress_address_offset[0] (
	.dataa(!\Add2~13_sumout ),
	.datab(!mem_81_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_burst_uncompress_address_offset[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_burst_uncompress_address_offset[0] .extended_lut = "off";
defparam \p1_burst_uncompress_address_offset[0] .lut_mask = 64'h1111111111111111;
defparam \p1_burst_uncompress_address_offset[0] .shared_arith = "off";

dffeas \burst_uncompress_address_offset[0] (
	.clk(clk),
	.d(\p1_burst_uncompress_address_offset[0]~combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sink_ready~0_combout ),
	.q(\burst_uncompress_address_offset[0]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_offset[0] .is_wysiwyg = "true";
defparam \burst_uncompress_address_offset[0] .power_up = "low";

cyclonev_lcell_comb \Add2~9 (
	.dataa(!comb),
	.datab(!burst_uncompress_busy1),
	.datac(!mem_37_0),
	.datad(!\Decoder0~2_combout ),
	.datae(gnd),
	.dataf(!\burst_uncompress_address_offset[1]~q ),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h0000FB40000000FF;
defparam \Add2~9 .shared_arith = "off";

cyclonev_lcell_comb \p1_burst_uncompress_address_offset[1] (
	.dataa(!\Add2~9_sumout ),
	.datab(!mem_82_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_burst_uncompress_address_offset[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_burst_uncompress_address_offset[1] .extended_lut = "off";
defparam \p1_burst_uncompress_address_offset[1] .lut_mask = 64'h1111111111111111;
defparam \p1_burst_uncompress_address_offset[1] .shared_arith = "off";

dffeas \burst_uncompress_address_offset[1] (
	.clk(clk),
	.d(\p1_burst_uncompress_address_offset[1]~combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sink_ready~0_combout ),
	.q(\burst_uncompress_address_offset[1]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_offset[1] .is_wysiwyg = "true";
defparam \burst_uncompress_address_offset[1] .power_up = "low";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!comb),
	.datab(!burst_uncompress_busy1),
	.datac(!mem_38_0),
	.datad(!\Decoder0~0_combout ),
	.datae(gnd),
	.dataf(!\burst_uncompress_address_offset[2]~q ),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h0000FB40000000FF;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \p1_burst_uncompress_address_offset[2] (
	.dataa(!mem_83_0),
	.datab(!\Add2~1_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_burst_uncompress_address_offset[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_burst_uncompress_address_offset[2] .extended_lut = "off";
defparam \p1_burst_uncompress_address_offset[2] .lut_mask = 64'h1111111111111111;
defparam \p1_burst_uncompress_address_offset[2] .shared_arith = "off";

dffeas \burst_uncompress_address_offset[2] (
	.clk(clk),
	.d(\p1_burst_uncompress_address_offset[2]~combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sink_ready~0_combout ),
	.q(\burst_uncompress_address_offset[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_offset[2] .is_wysiwyg = "true";
defparam \burst_uncompress_address_offset[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_address_base~1 (
	.dataa(!mem_39_0),
	.datab(!mem_84_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_address_base~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_address_base~1 .extended_lut = "off";
defparam \burst_uncompress_address_base~1 .lut_mask = 64'h4444444444444444;
defparam \burst_uncompress_address_base~1 .shared_arith = "off";

dffeas \burst_uncompress_address_base[3] (
	.clk(clk),
	.d(\burst_uncompress_address_base~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\burst_uncompress_address_base[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_base[3] .is_wysiwyg = "true";
defparam \burst_uncompress_address_base[3] .power_up = "low";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!mem_90_0),
	.datab(!mem_91_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'h1111111111111111;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add2~5 (
	.dataa(!comb),
	.datab(!burst_uncompress_busy1),
	.datac(!mem_39_0),
	.datad(!\Decoder0~1_combout ),
	.datae(gnd),
	.dataf(!\burst_uncompress_address_offset[3]~q ),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h0000FB40000000FF;
defparam \Add2~5 .shared_arith = "off";

cyclonev_lcell_comb \p1_burst_uncompress_address_offset[3] (
	.dataa(!mem_84_0),
	.datab(!\Add2~5_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p1_burst_uncompress_address_offset[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_burst_uncompress_address_offset[3] .extended_lut = "off";
defparam \p1_burst_uncompress_address_offset[3] .lut_mask = 64'h1111111111111111;
defparam \p1_burst_uncompress_address_offset[3] .shared_arith = "off";

dffeas \burst_uncompress_address_offset[3] (
	.clk(clk),
	.d(\p1_burst_uncompress_address_offset[3]~combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sink_ready~0_combout ),
	.q(\burst_uncompress_address_offset[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_address_offset[3] .is_wysiwyg = "true";
defparam \burst_uncompress_address_offset[3] .power_up = "low";

endmodule

module Computer_System_altera_merlin_slave_translator_1 (
	clk,
	in_ready_hold,
	mem_used_1,
	out_valid_reg,
	read_latency_shift_reg_0,
	reset,
	in_data_reg_69,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	in_ready_hold;
input 	mem_used_1;
input 	out_valid_reg;
output 	read_latency_shift_reg_0;
input 	reset;
input 	in_data_reg_69;
input 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!in_ready_hold),
	.datab(!out_valid_reg),
	.datac(!WideOr0),
	.datad(!mem_used_1),
	.datae(!in_data_reg_69),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0000100000001000;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_traffic_limiter (
	h2f_ARVALID_0,
	h2f_RREADY_0,
	clk,
	saved_grant_1,
	in_ready,
	sink1_ready,
	nxt_in_ready,
	out_valid,
	src_payload,
	src0_valid,
	src_payload_0,
	WideOr1,
	cmd_src_valid_1,
	reset,
	src_payload1)/* synthesis synthesis_greybox=0 */;
input 	h2f_ARVALID_0;
input 	h2f_RREADY_0;
input 	clk;
input 	saved_grant_1;
input 	in_ready;
input 	sink1_ready;
input 	nxt_in_ready;
input 	out_valid;
input 	src_payload;
input 	src0_valid;
input 	src_payload_0;
input 	WideOr1;
output 	cmd_src_valid_1;
input 	reset;
input 	src_payload1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \last_channel[1]~0_combout ;
wire \last_channel[1]~q ;
wire \pending_response_count[0]~1_combout ;
wire \response_sink_accepted~0_combout ;
wire \pending_response_count[1]~0_combout ;
wire \pending_response_count[0]~q ;
wire \Add0~0_combout ;
wire \pending_response_count[1]~q ;
wire \response_sink_accepted~combout ;
wire \has_pending_responses~0_combout ;
wire \has_pending_responses~q ;


cyclonev_lcell_comb \cmd_src_valid[1]~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!\last_channel[1]~q ),
	.datac(!\has_pending_responses~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cmd_src_valid_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_src_valid[1]~0 .extended_lut = "off";
defparam \cmd_src_valid[1]~0 .lut_mask = 64'h5151515151515151;
defparam \cmd_src_valid[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \last_channel[1]~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!\last_channel[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_channel[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_channel[1]~0 .extended_lut = "off";
defparam \last_channel[1]~0 .lut_mask = 64'h7777777777777777;
defparam \last_channel[1]~0 .shared_arith = "off";

dffeas \last_channel[1] (
	.clk(clk),
	.d(\last_channel[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_channel[1]~q ),
	.prn(vcc));
defparam \last_channel[1] .is_wysiwyg = "true";
defparam \last_channel[1] .power_up = "low";

cyclonev_lcell_comb \pending_response_count[0]~1 (
	.dataa(!\pending_response_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~1 .extended_lut = "off";
defparam \pending_response_count[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \pending_response_count[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~0 (
	.dataa(!h2f_RREADY_0),
	.datab(!out_valid),
	.datac(!src_payload),
	.datad(gnd),
	.datae(!src0_valid),
	.dataf(!src_payload1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~0 .extended_lut = "off";
defparam \response_sink_accepted~0 .lut_mask = 64'h0404000055555555;
defparam \response_sink_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[1]~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!saved_grant_1),
	.datac(!in_ready),
	.datad(!nxt_in_ready),
	.datae(!WideOr1),
	.dataf(!\response_sink_accepted~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[1]~0 .extended_lut = "off";
defparam \pending_response_count[1]~0 .lut_mask = 64'h100010001000EFFF;
defparam \pending_response_count[1]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!WideOr1),
	.datab(!\pending_response_count[1]~q ),
	.datac(!\pending_response_count[0]~q ),
	.datad(!\response_sink_accepted~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h3C693C693C693C69;
defparam \Add0~0 .shared_arith = "off";

dffeas \pending_response_count[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[1]~q ),
	.prn(vcc));
defparam \pending_response_count[1] .is_wysiwyg = "true";
defparam \pending_response_count[1] .power_up = "low";

cyclonev_lcell_comb response_sink_accepted(
	.dataa(!h2f_RREADY_0),
	.datab(!src_payload_0),
	.datac(!WideOr1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam response_sink_accepted.extended_lut = "off";
defparam response_sink_accepted.lut_mask = 64'h0101010101010101;
defparam response_sink_accepted.shared_arith = "off";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!h2f_ARVALID_0),
	.datab(!sink1_ready),
	.datac(!\has_pending_responses~q ),
	.datad(!\pending_response_count[1]~q ),
	.datae(!\pending_response_count[0]~q ),
	.dataf(!\response_sink_accepted~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'h1F0F0F0F0F0F010F;
defparam \has_pending_responses~0 .shared_arith = "off";

dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\has_pending_responses~q ),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

endmodule

module Computer_System_altera_merlin_traffic_limiter_1 (
	h2f_BREADY_0,
	h2f_WLAST_0,
	clk,
	Equal0,
	Equal01,
	Equal02,
	sink_ready,
	last_channel_0,
	has_pending_responses1,
	cmd_sink_ready,
	out_valid,
	src_payload,
	src0_valid,
	mem_126_0,
	src0_valid1,
	WideOr1,
	last_cycle,
	cmd_sink_channel,
	last_channel_1,
	reset,
	sink_ready1)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_WLAST_0;
input 	clk;
input 	Equal0;
input 	Equal01;
input 	Equal02;
input 	sink_ready;
output 	last_channel_0;
output 	has_pending_responses1;
output 	cmd_sink_ready;
input 	out_valid;
input 	src_payload;
input 	src0_valid;
input 	mem_126_0;
input 	src0_valid1;
input 	WideOr1;
input 	last_cycle;
input 	[1:0] cmd_sink_channel;
output 	last_channel_1;
input 	reset;
input 	sink_ready1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \save_dest_id~0_combout ;
wire \pending_response_count[0]~1_combout ;
wire \response_sink_accepted~0_combout ;
wire \response_sink_accepted~1_combout ;
wire \pending_response_count[1]~0_combout ;
wire \pending_response_count[0]~q ;
wire \Add0~0_combout ;
wire \pending_response_count[1]~q ;
wire \has_pending_responses~0_combout ;
wire \has_pending_responses~1_combout ;
wire \has_pending_responses~2_combout ;
wire \last_channel[1]~0_combout ;


dffeas \last_channel[0] (
	.clk(clk),
	.d(cmd_sink_channel[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_0),
	.prn(vcc));
defparam \last_channel[0] .is_wysiwyg = "true";
defparam \last_channel[0] .power_up = "low";

dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

cyclonev_lcell_comb \cmd_sink_ready~0 (
	.dataa(!Equal0),
	.datab(!Equal01),
	.datac(!Equal02),
	.datad(!last_channel_0),
	.datae(!has_pending_responses1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cmd_sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_sink_ready~0 .extended_lut = "off";
defparam \cmd_sink_ready~0 .lut_mask = 64'h000001FE000001FE;
defparam \cmd_sink_ready~0 .shared_arith = "off";

dffeas \last_channel[1] (
	.clk(clk),
	.d(\last_channel[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_1),
	.prn(vcc));
defparam \last_channel[1] .is_wysiwyg = "true";
defparam \last_channel[1] .power_up = "low";

cyclonev_lcell_comb \save_dest_id~0 (
	.dataa(!Equal0),
	.datab(!Equal01),
	.datac(!Equal02),
	.datad(!last_channel_0),
	.datae(!has_pending_responses1),
	.dataf(!last_cycle),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\save_dest_id~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \save_dest_id~0 .extended_lut = "off";
defparam \save_dest_id~0 .lut_mask = 64'h00000000FFFFFE01;
defparam \save_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[0]~1 (
	.dataa(!\pending_response_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~1 .extended_lut = "off";
defparam \pending_response_count[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \pending_response_count[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~0 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(gnd),
	.datad(!src0_valid),
	.datae(!mem_126_0),
	.dataf(!src0_valid1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~0 .extended_lut = "off";
defparam \response_sink_accepted~0 .lut_mask = 64'h002200220022FFFF;
defparam \response_sink_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~1 (
	.dataa(!h2f_BREADY_0),
	.datab(!WideOr1),
	.datac(!\response_sink_accepted~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~1 .extended_lut = "off";
defparam \response_sink_accepted~1 .lut_mask = 64'h0101010101010101;
defparam \response_sink_accepted~1 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[1]~0 (
	.dataa(!h2f_WLAST_0),
	.datab(!sink_ready1),
	.datac(!sink_ready),
	.datad(!\save_dest_id~0_combout ),
	.datae(!\response_sink_accepted~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[1]~0 .extended_lut = "off";
defparam \pending_response_count[1]~0 .lut_mask = 64'h0015FFEA0015FFEA;
defparam \pending_response_count[1]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!WideOr1),
	.datac(!\pending_response_count[1]~q ),
	.datad(!\pending_response_count[0]~q ),
	.datae(!\response_sink_accepted~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h0FF01EE10FF01EE1;
defparam \Add0~0 .shared_arith = "off";

dffeas \pending_response_count[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[1]~q ),
	.prn(vcc));
defparam \pending_response_count[1] .is_wysiwyg = "true";
defparam \pending_response_count[1] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!has_pending_responses1),
	.datac(!WideOr1),
	.datad(!\pending_response_count[1]~q ),
	.datae(!\pending_response_count[0]~q ),
	.dataf(!\response_sink_accepted~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'h3333333333333233;
defparam \has_pending_responses~0 .shared_arith = "off";

cyclonev_lcell_comb \has_pending_responses~1 (
	.dataa(!h2f_BREADY_0),
	.datab(!has_pending_responses1),
	.datac(!WideOr1),
	.datad(!\pending_response_count[1]~q ),
	.datae(!\pending_response_count[0]~q ),
	.dataf(!\response_sink_accepted~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~1 .extended_lut = "off";
defparam \has_pending_responses~1 .lut_mask = 64'h00CCCCCC04CCCCCC;
defparam \has_pending_responses~1 .shared_arith = "off";

cyclonev_lcell_comb \has_pending_responses~2 (
	.dataa(!h2f_WLAST_0),
	.datab(!sink_ready1),
	.datac(!sink_ready),
	.datad(!\save_dest_id~0_combout ),
	.datae(!\has_pending_responses~0_combout ),
	.dataf(!\has_pending_responses~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~2 .extended_lut = "off";
defparam \has_pending_responses~2 .lut_mask = 64'h0015FFFF0000FFFF;
defparam \has_pending_responses~2 .shared_arith = "off";

cyclonev_lcell_comb \last_channel[1]~0 (
	.dataa(!cmd_sink_channel[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_channel[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_channel[1]~0 .extended_lut = "off";
defparam \last_channel[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \last_channel[1]~0 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_width_adapter (
	h2f_WLAST_0,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WDATA_1,
	h2f_WDATA_2,
	h2f_WDATA_3,
	h2f_WDATA_4,
	h2f_WDATA_5,
	h2f_WDATA_6,
	h2f_WDATA_7,
	h2f_WDATA_8,
	h2f_WDATA_9,
	h2f_WDATA_10,
	h2f_WDATA_11,
	h2f_WDATA_12,
	h2f_WDATA_13,
	h2f_WDATA_14,
	h2f_WDATA_15,
	h2f_WDATA_16,
	h2f_WDATA_17,
	h2f_WDATA_18,
	h2f_WDATA_19,
	h2f_WDATA_20,
	h2f_WDATA_21,
	h2f_WDATA_22,
	h2f_WDATA_23,
	h2f_WDATA_24,
	h2f_WDATA_25,
	h2f_WDATA_26,
	h2f_WDATA_27,
	h2f_WDATA_28,
	h2f_WDATA_29,
	h2f_WDATA_30,
	h2f_WDATA_31,
	h2f_WDATA_32,
	h2f_WDATA_33,
	h2f_WDATA_34,
	h2f_WDATA_35,
	h2f_WDATA_36,
	h2f_WDATA_37,
	h2f_WDATA_38,
	h2f_WDATA_39,
	h2f_WDATA_40,
	h2f_WDATA_41,
	h2f_WDATA_42,
	h2f_WDATA_43,
	h2f_WDATA_44,
	h2f_WDATA_45,
	h2f_WDATA_46,
	h2f_WDATA_47,
	h2f_WDATA_48,
	h2f_WDATA_49,
	h2f_WDATA_50,
	h2f_WDATA_51,
	h2f_WDATA_52,
	h2f_WDATA_53,
	h2f_WDATA_54,
	h2f_WDATA_55,
	h2f_WDATA_56,
	h2f_WDATA_57,
	h2f_WDATA_58,
	h2f_WDATA_59,
	h2f_WDATA_60,
	h2f_WDATA_61,
	h2f_WDATA_62,
	h2f_WDATA_63,
	h2f_WDATA_64,
	h2f_WDATA_65,
	h2f_WDATA_66,
	h2f_WDATA_67,
	h2f_WDATA_68,
	h2f_WDATA_69,
	h2f_WDATA_70,
	h2f_WDATA_71,
	h2f_WDATA_72,
	h2f_WDATA_73,
	h2f_WDATA_74,
	h2f_WDATA_75,
	h2f_WDATA_76,
	h2f_WDATA_77,
	h2f_WDATA_78,
	h2f_WDATA_79,
	h2f_WDATA_80,
	h2f_WDATA_81,
	h2f_WDATA_82,
	h2f_WDATA_83,
	h2f_WDATA_84,
	h2f_WDATA_85,
	h2f_WDATA_86,
	h2f_WDATA_87,
	h2f_WDATA_88,
	h2f_WDATA_89,
	h2f_WDATA_90,
	h2f_WDATA_91,
	h2f_WDATA_92,
	h2f_WDATA_93,
	h2f_WDATA_94,
	h2f_WDATA_95,
	h2f_WDATA_96,
	h2f_WDATA_97,
	h2f_WDATA_98,
	h2f_WDATA_99,
	h2f_WDATA_100,
	h2f_WDATA_101,
	h2f_WDATA_102,
	h2f_WDATA_103,
	h2f_WDATA_104,
	h2f_WDATA_105,
	h2f_WDATA_106,
	h2f_WDATA_107,
	h2f_WDATA_108,
	h2f_WDATA_109,
	h2f_WDATA_110,
	h2f_WDATA_111,
	h2f_WDATA_112,
	h2f_WDATA_113,
	h2f_WDATA_114,
	h2f_WDATA_115,
	h2f_WDATA_116,
	h2f_WDATA_117,
	h2f_WDATA_118,
	h2f_WDATA_119,
	h2f_WDATA_120,
	h2f_WDATA_121,
	h2f_WDATA_122,
	h2f_WDATA_123,
	h2f_WDATA_124,
	h2f_WDATA_125,
	h2f_WDATA_126,
	h2f_WDATA_127,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	h2f_WSTRB_4,
	h2f_WSTRB_5,
	h2f_WSTRB_6,
	h2f_WSTRB_7,
	h2f_WSTRB_8,
	h2f_WSTRB_9,
	h2f_WSTRB_10,
	h2f_WSTRB_11,
	h2f_WSTRB_12,
	h2f_WSTRB_13,
	h2f_WSTRB_14,
	h2f_WSTRB_15,
	outclk_wire_0,
	out_data_37,
	Mux4,
	Mux5,
	Mux6,
	Mux7,
	Mux8,
	Mux9,
	Mux10,
	Mux11,
	Mux12,
	Mux13,
	Mux14,
	Mux15,
	Mux16,
	Mux17,
	Mux18,
	Mux19,
	Mux20,
	Mux21,
	Mux22,
	Mux23,
	Mux24,
	Mux25,
	Mux26,
	Mux27,
	Mux28,
	Mux29,
	Mux30,
	Mux31,
	Mux32,
	Mux33,
	Mux34,
	Mux35,
	Mux3,
	Mux2,
	Mux1,
	Mux0,
	in_ready_hold,
	Equal0,
	Equal01,
	Equal02,
	nxt_in_ready,
	out_valid_reg,
	saved_grant_0,
	count_1,
	count_0,
	r_sync_rst,
	out_data_2,
	out_data_3,
	src0_valid,
	LessThan2,
	int_output_sel_0,
	int_output_sel_1,
	src_payload,
	src_payload1,
	src_payload2,
	cp_ready,
	out_data_1,
	Decoder0,
	out_data_0,
	out_endofpacket,
	nxt_in_ready1,
	nxt_in_ready2,
	src0_valid1,
	out_data_90,
	out_data_91,
	out_data_36)/* synthesis synthesis_greybox=0 */;
input 	h2f_WLAST_0;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WDATA_1;
input 	h2f_WDATA_2;
input 	h2f_WDATA_3;
input 	h2f_WDATA_4;
input 	h2f_WDATA_5;
input 	h2f_WDATA_6;
input 	h2f_WDATA_7;
input 	h2f_WDATA_8;
input 	h2f_WDATA_9;
input 	h2f_WDATA_10;
input 	h2f_WDATA_11;
input 	h2f_WDATA_12;
input 	h2f_WDATA_13;
input 	h2f_WDATA_14;
input 	h2f_WDATA_15;
input 	h2f_WDATA_16;
input 	h2f_WDATA_17;
input 	h2f_WDATA_18;
input 	h2f_WDATA_19;
input 	h2f_WDATA_20;
input 	h2f_WDATA_21;
input 	h2f_WDATA_22;
input 	h2f_WDATA_23;
input 	h2f_WDATA_24;
input 	h2f_WDATA_25;
input 	h2f_WDATA_26;
input 	h2f_WDATA_27;
input 	h2f_WDATA_28;
input 	h2f_WDATA_29;
input 	h2f_WDATA_30;
input 	h2f_WDATA_31;
input 	h2f_WDATA_32;
input 	h2f_WDATA_33;
input 	h2f_WDATA_34;
input 	h2f_WDATA_35;
input 	h2f_WDATA_36;
input 	h2f_WDATA_37;
input 	h2f_WDATA_38;
input 	h2f_WDATA_39;
input 	h2f_WDATA_40;
input 	h2f_WDATA_41;
input 	h2f_WDATA_42;
input 	h2f_WDATA_43;
input 	h2f_WDATA_44;
input 	h2f_WDATA_45;
input 	h2f_WDATA_46;
input 	h2f_WDATA_47;
input 	h2f_WDATA_48;
input 	h2f_WDATA_49;
input 	h2f_WDATA_50;
input 	h2f_WDATA_51;
input 	h2f_WDATA_52;
input 	h2f_WDATA_53;
input 	h2f_WDATA_54;
input 	h2f_WDATA_55;
input 	h2f_WDATA_56;
input 	h2f_WDATA_57;
input 	h2f_WDATA_58;
input 	h2f_WDATA_59;
input 	h2f_WDATA_60;
input 	h2f_WDATA_61;
input 	h2f_WDATA_62;
input 	h2f_WDATA_63;
input 	h2f_WDATA_64;
input 	h2f_WDATA_65;
input 	h2f_WDATA_66;
input 	h2f_WDATA_67;
input 	h2f_WDATA_68;
input 	h2f_WDATA_69;
input 	h2f_WDATA_70;
input 	h2f_WDATA_71;
input 	h2f_WDATA_72;
input 	h2f_WDATA_73;
input 	h2f_WDATA_74;
input 	h2f_WDATA_75;
input 	h2f_WDATA_76;
input 	h2f_WDATA_77;
input 	h2f_WDATA_78;
input 	h2f_WDATA_79;
input 	h2f_WDATA_80;
input 	h2f_WDATA_81;
input 	h2f_WDATA_82;
input 	h2f_WDATA_83;
input 	h2f_WDATA_84;
input 	h2f_WDATA_85;
input 	h2f_WDATA_86;
input 	h2f_WDATA_87;
input 	h2f_WDATA_88;
input 	h2f_WDATA_89;
input 	h2f_WDATA_90;
input 	h2f_WDATA_91;
input 	h2f_WDATA_92;
input 	h2f_WDATA_93;
input 	h2f_WDATA_94;
input 	h2f_WDATA_95;
input 	h2f_WDATA_96;
input 	h2f_WDATA_97;
input 	h2f_WDATA_98;
input 	h2f_WDATA_99;
input 	h2f_WDATA_100;
input 	h2f_WDATA_101;
input 	h2f_WDATA_102;
input 	h2f_WDATA_103;
input 	h2f_WDATA_104;
input 	h2f_WDATA_105;
input 	h2f_WDATA_106;
input 	h2f_WDATA_107;
input 	h2f_WDATA_108;
input 	h2f_WDATA_109;
input 	h2f_WDATA_110;
input 	h2f_WDATA_111;
input 	h2f_WDATA_112;
input 	h2f_WDATA_113;
input 	h2f_WDATA_114;
input 	h2f_WDATA_115;
input 	h2f_WDATA_116;
input 	h2f_WDATA_117;
input 	h2f_WDATA_118;
input 	h2f_WDATA_119;
input 	h2f_WDATA_120;
input 	h2f_WDATA_121;
input 	h2f_WDATA_122;
input 	h2f_WDATA_123;
input 	h2f_WDATA_124;
input 	h2f_WDATA_125;
input 	h2f_WDATA_126;
input 	h2f_WDATA_127;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
input 	h2f_WSTRB_4;
input 	h2f_WSTRB_5;
input 	h2f_WSTRB_6;
input 	h2f_WSTRB_7;
input 	h2f_WSTRB_8;
input 	h2f_WSTRB_9;
input 	h2f_WSTRB_10;
input 	h2f_WSTRB_11;
input 	h2f_WSTRB_12;
input 	h2f_WSTRB_13;
input 	h2f_WSTRB_14;
input 	h2f_WSTRB_15;
input 	outclk_wire_0;
output 	out_data_37;
output 	Mux4;
output 	Mux5;
output 	Mux6;
output 	Mux7;
output 	Mux8;
output 	Mux9;
output 	Mux10;
output 	Mux11;
output 	Mux12;
output 	Mux13;
output 	Mux14;
output 	Mux15;
output 	Mux16;
output 	Mux17;
output 	Mux18;
output 	Mux19;
output 	Mux20;
output 	Mux21;
output 	Mux22;
output 	Mux23;
output 	Mux24;
output 	Mux25;
output 	Mux26;
output 	Mux27;
output 	Mux28;
output 	Mux29;
output 	Mux30;
output 	Mux31;
output 	Mux32;
output 	Mux33;
output 	Mux34;
output 	Mux35;
output 	Mux3;
output 	Mux2;
output 	Mux1;
output 	Mux0;
input 	in_ready_hold;
input 	Equal0;
input 	Equal01;
input 	Equal02;
input 	nxt_in_ready;
input 	out_valid_reg;
input 	saved_grant_0;
output 	count_1;
output 	count_0;
input 	r_sync_rst;
input 	out_data_2;
input 	out_data_3;
input 	src0_valid;
input 	LessThan2;
output 	int_output_sel_0;
output 	int_output_sel_1;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	cp_ready;
input 	out_data_1;
input 	Decoder0;
input 	out_data_0;
output 	out_endofpacket;
input 	nxt_in_ready1;
input 	nxt_in_ready2;
input 	src0_valid1;
output 	out_data_90;
output 	out_data_91;
output 	out_data_36;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Decoder0~2_combout ;
wire \Decoder0~3_combout ;
wire \LessThan3~0_combout ;
wire \Decoder0~4_combout ;
wire \Add1~14 ;
wire \Add1~9_sumout ;
wire \out_endofpacket~0_combout ;
wire \use_reg~0_combout ;
wire \use_reg~q ;
wire \address_reg~0_combout ;
wire \address_reg[1]~q ;
wire \Decoder0~0_combout ;
wire \Decoder0~1_combout ;
wire \Add0~0_combout ;
wire \Add0~1_combout ;
wire \count~0_combout ;
wire \count~1_combout ;
wire \Add1~10 ;
wire \Add1~1_sumout ;
wire \address_reg[2]~q ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \address_reg[3]~q ;
wire \endofpacket_reg~0_combout ;
wire \endofpacket_reg~q ;
wire \Add1~13_sumout ;
wire \address_reg[0]~q ;


cyclonev_lcell_comb \out_data[37]~3 (
	.dataa(!h2f_AWSIZE_2),
	.datab(!h2f_AWSIZE_1),
	.datac(!\address_reg[1]~q ),
	.datad(!h2f_AWSIZE_0),
	.datae(!\use_reg~q ),
	.dataf(!saved_grant_0),
	.datag(!out_data_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_37),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[37]~3 .extended_lut = "on";
defparam \out_data[37]~3 .lut_mask = 64'h00000F0F0A080F0F;
defparam \out_data[37]~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux4~0 (
	.dataa(!h2f_WDATA_127),
	.datab(!h2f_WDATA_63),
	.datac(!h2f_WDATA_95),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_31),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~0 .extended_lut = "on";
defparam \Mux4~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux4~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux5~0 (
	.dataa(!h2f_WDATA_126),
	.datab(!h2f_WDATA_62),
	.datac(!h2f_WDATA_94),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_30),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux5),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~0 .extended_lut = "on";
defparam \Mux5~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux5~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux6~0 (
	.dataa(!h2f_WDATA_125),
	.datab(!h2f_WDATA_61),
	.datac(!h2f_WDATA_93),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_29),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux6),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~0 .extended_lut = "on";
defparam \Mux6~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux6~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux7~0 (
	.dataa(!h2f_WDATA_124),
	.datab(!h2f_WDATA_60),
	.datac(!h2f_WDATA_92),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_28),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux7),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~0 .extended_lut = "on";
defparam \Mux7~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux7~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~0 (
	.dataa(!h2f_WDATA_123),
	.datab(!h2f_WDATA_59),
	.datac(!h2f_WDATA_91),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_27),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux8),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~0 .extended_lut = "on";
defparam \Mux8~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux8~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux9~0 (
	.dataa(!h2f_WDATA_122),
	.datab(!h2f_WDATA_58),
	.datac(!h2f_WDATA_90),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_26),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux9),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~0 .extended_lut = "on";
defparam \Mux9~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux9~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux10~0 (
	.dataa(!h2f_WDATA_121),
	.datab(!h2f_WDATA_57),
	.datac(!h2f_WDATA_89),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_25),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux10),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~0 .extended_lut = "on";
defparam \Mux10~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux10~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux11~0 (
	.dataa(!h2f_WDATA_120),
	.datab(!h2f_WDATA_56),
	.datac(!h2f_WDATA_88),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_24),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~0 .extended_lut = "on";
defparam \Mux11~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux11~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux12~0 (
	.dataa(!h2f_WDATA_119),
	.datab(!h2f_WDATA_55),
	.datac(!h2f_WDATA_87),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_23),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux12),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux12~0 .extended_lut = "on";
defparam \Mux12~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux12~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux13~0 (
	.dataa(!h2f_WDATA_118),
	.datab(!h2f_WDATA_54),
	.datac(!h2f_WDATA_86),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_22),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux13),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~0 .extended_lut = "on";
defparam \Mux13~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux13~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux14~0 (
	.dataa(!h2f_WDATA_117),
	.datab(!h2f_WDATA_53),
	.datac(!h2f_WDATA_85),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_21),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux14),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~0 .extended_lut = "on";
defparam \Mux14~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux14~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux15~0 (
	.dataa(!h2f_WDATA_116),
	.datab(!h2f_WDATA_52),
	.datac(!h2f_WDATA_84),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_20),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux15),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux15~0 .extended_lut = "on";
defparam \Mux15~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux15~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux16~0 (
	.dataa(!h2f_WDATA_115),
	.datab(!h2f_WDATA_51),
	.datac(!h2f_WDATA_83),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_19),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux16),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~0 .extended_lut = "on";
defparam \Mux16~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux16~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux17~0 (
	.dataa(!h2f_WDATA_114),
	.datab(!h2f_WDATA_50),
	.datac(!h2f_WDATA_82),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_18),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux17),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux17~0 .extended_lut = "on";
defparam \Mux17~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux17~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux18~0 (
	.dataa(!h2f_WDATA_113),
	.datab(!h2f_WDATA_49),
	.datac(!h2f_WDATA_81),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_17),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux18),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux18~0 .extended_lut = "on";
defparam \Mux18~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux18~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux19~0 (
	.dataa(!h2f_WDATA_112),
	.datab(!h2f_WDATA_48),
	.datac(!h2f_WDATA_80),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_16),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux19),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux19~0 .extended_lut = "on";
defparam \Mux19~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux19~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux20~0 (
	.dataa(!h2f_WDATA_111),
	.datab(!h2f_WDATA_47),
	.datac(!h2f_WDATA_79),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_15),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux20),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux20~0 .extended_lut = "on";
defparam \Mux20~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux20~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux21~0 (
	.dataa(!h2f_WDATA_110),
	.datab(!h2f_WDATA_46),
	.datac(!h2f_WDATA_78),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_14),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux21),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux21~0 .extended_lut = "on";
defparam \Mux21~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux21~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux22~0 (
	.dataa(!h2f_WDATA_109),
	.datab(!h2f_WDATA_45),
	.datac(!h2f_WDATA_77),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_13),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux22),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~0 .extended_lut = "on";
defparam \Mux22~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux22~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux23~0 (
	.dataa(!h2f_WDATA_108),
	.datab(!h2f_WDATA_44),
	.datac(!h2f_WDATA_76),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_12),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux23),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux23~0 .extended_lut = "on";
defparam \Mux23~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux23~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~0 (
	.dataa(!h2f_WDATA_107),
	.datab(!h2f_WDATA_43),
	.datac(!h2f_WDATA_75),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_11),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux24),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~0 .extended_lut = "on";
defparam \Mux24~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux24~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux25~0 (
	.dataa(!h2f_WDATA_106),
	.datab(!h2f_WDATA_42),
	.datac(!h2f_WDATA_74),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_10),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux25),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~0 .extended_lut = "on";
defparam \Mux25~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux25~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux26~0 (
	.dataa(!h2f_WDATA_105),
	.datab(!h2f_WDATA_41),
	.datac(!h2f_WDATA_73),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_9),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux26),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~0 .extended_lut = "on";
defparam \Mux26~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux26~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux27~0 (
	.dataa(!h2f_WDATA_104),
	.datab(!h2f_WDATA_40),
	.datac(!h2f_WDATA_72),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_8),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux27),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~0 .extended_lut = "on";
defparam \Mux27~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux27~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux28~0 (
	.dataa(!h2f_WDATA_103),
	.datab(!h2f_WDATA_39),
	.datac(!h2f_WDATA_71),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_7),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux28),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux28~0 .extended_lut = "on";
defparam \Mux28~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux28~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux29~0 (
	.dataa(!h2f_WDATA_102),
	.datab(!h2f_WDATA_38),
	.datac(!h2f_WDATA_70),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_6),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux29),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux29~0 .extended_lut = "on";
defparam \Mux29~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux29~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux30~0 (
	.dataa(!h2f_WDATA_101),
	.datab(!h2f_WDATA_37),
	.datac(!h2f_WDATA_69),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_5),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux30),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux30~0 .extended_lut = "on";
defparam \Mux30~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux30~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux31~0 (
	.dataa(!h2f_WDATA_100),
	.datab(!h2f_WDATA_36),
	.datac(!h2f_WDATA_68),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_4),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux31),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux31~0 .extended_lut = "on";
defparam \Mux31~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux31~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~0 (
	.dataa(!h2f_WDATA_99),
	.datab(!h2f_WDATA_35),
	.datac(!h2f_WDATA_67),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_3),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux32),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~0 .extended_lut = "on";
defparam \Mux32~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux32~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux33~0 (
	.dataa(!h2f_WDATA_98),
	.datab(!h2f_WDATA_34),
	.datac(!h2f_WDATA_66),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_2),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux33),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux33~0 .extended_lut = "on";
defparam \Mux33~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux33~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux34~0 (
	.dataa(!h2f_WDATA_97),
	.datab(!h2f_WDATA_33),
	.datac(!h2f_WDATA_65),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux34),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux34~0 .extended_lut = "on";
defparam \Mux34~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux34~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux35~0 (
	.dataa(!h2f_WDATA_96),
	.datab(!h2f_WDATA_32),
	.datac(!h2f_WDATA_64),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_0),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux35),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux35~0 .extended_lut = "on";
defparam \Mux35~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux35~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~0 (
	.dataa(!h2f_WSTRB_12),
	.datab(!h2f_WSTRB_4),
	.datac(!h2f_WSTRB_8),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WSTRB_0),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "on";
defparam \Mux3~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux3~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~0 (
	.dataa(!h2f_WSTRB_13),
	.datab(!h2f_WSTRB_5),
	.datac(!h2f_WSTRB_9),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WSTRB_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~0 .extended_lut = "on";
defparam \Mux2~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux2~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux1~0 (
	.dataa(!h2f_WSTRB_14),
	.datab(!h2f_WSTRB_6),
	.datac(!h2f_WSTRB_10),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WSTRB_2),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~0 .extended_lut = "on";
defparam \Mux1~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux1~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!h2f_WSTRB_15),
	.datab(!h2f_WSTRB_7),
	.datac(!h2f_WSTRB_11),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WSTRB_3),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "on";
defparam \Mux0~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux0~0 .shared_arith = "off";

dffeas \count[1] (
	.clk(outclk_wire_0),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count~1_combout ),
	.q(count_1),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

dffeas \count[0] (
	.clk(outclk_wire_0),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count~1_combout ),
	.q(count_0),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cyclonev_lcell_comb \int_output_sel[0]~0 (
	.dataa(!out_data_2),
	.datab(!saved_grant_0),
	.datac(!LessThan2),
	.datad(!\address_reg[2]~q ),
	.datae(!\use_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(int_output_sel_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_output_sel[0]~0 .extended_lut = "off";
defparam \int_output_sel[0]~0 .lut_mask = 64'h101000FF101000FF;
defparam \int_output_sel[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \int_output_sel[1]~1 (
	.dataa(!h2f_AWSIZE_2),
	.datab(!out_data_3),
	.datac(!saved_grant_0),
	.datad(!\use_reg~q ),
	.datae(!\address_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(int_output_sel_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_output_sel[1]~1 .extended_lut = "off";
defparam \int_output_sel[1]~1 .lut_mask = 64'h020002FF020002FF;
defparam \int_output_sel[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_endofpacket~1 (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_0),
	.datac(!LessThan2),
	.datad(!\out_endofpacket~0_combout ),
	.datae(!\use_reg~q ),
	.dataf(!\endofpacket_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_endofpacket),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_endofpacket~1 .extended_lut = "off";
defparam \out_endofpacket~1 .lut_mask = 64'h10101000101010FF;
defparam \out_endofpacket~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[90]~0 (
	.dataa(!src_payload),
	.datab(!src_payload1),
	.datac(!src_payload2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_90),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[90]~0 .extended_lut = "off";
defparam \out_data[90]~0 .lut_mask = 64'h2020202020202020;
defparam \out_data[90]~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[91]~1 (
	.dataa(!h2f_AWSIZE_1),
	.datab(!h2f_AWSIZE_2),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_91),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[91]~1 .extended_lut = "off";
defparam \out_data[91]~1 .lut_mask = 64'h0707070707070707;
defparam \out_data[91]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[36]~2 (
	.dataa(!saved_grant_0),
	.datab(!LessThan2),
	.datac(!Decoder0),
	.datad(!out_data_0),
	.datae(!\use_reg~q ),
	.dataf(!\address_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_36),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[36]~2 .extended_lut = "off";
defparam \out_data[36]~2 .lut_mask = 64'h004500000045FFFF;
defparam \out_data[36]~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~2 (
	.dataa(!src_payload),
	.datab(!src_payload1),
	.datac(!src_payload2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~2 .extended_lut = "off";
defparam \Decoder0~2 .lut_mask = 64'h0404040404040404;
defparam \Decoder0~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~3 (
	.dataa(!src_payload),
	.datab(!src_payload1),
	.datac(!src_payload2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~3 .extended_lut = "off";
defparam \Decoder0~3 .lut_mask = 64'h0101010101010101;
defparam \Decoder0~3 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~0 (
	.dataa(!src_payload),
	.datab(!src_payload2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~0 .extended_lut = "off";
defparam \LessThan3~0 .lut_mask = 64'h6666666666666666;
defparam \LessThan3~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~4 (
	.dataa(!src_payload),
	.datab(!src_payload1),
	.datac(!src_payload2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~4 .extended_lut = "off";
defparam \Decoder0~4 .lut_mask = 64'h8080808080808080;
defparam \Decoder0~4 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(!\Decoder0~2_combout ),
	.datab(!\Decoder0~3_combout ),
	.datac(!\Decoder0~4_combout ),
	.datad(!out_data_36),
	.datae(gnd),
	.dataf(!\LessThan3~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000F7FF000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(!\Decoder0~2_combout ),
	.datab(!\Decoder0~3_combout ),
	.datac(!out_data_90),
	.datad(!out_data_37),
	.datae(gnd),
	.dataf(!\LessThan3~0_combout ),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000F7FF000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \out_endofpacket~0 (
	.dataa(!count_1),
	.datab(!count_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_endofpacket~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_endofpacket~0 .extended_lut = "off";
defparam \out_endofpacket~0 .lut_mask = 64'h2222222222222222;
defparam \out_endofpacket~0 .shared_arith = "off";

cyclonev_lcell_comb \use_reg~0 (
	.dataa(!LessThan2),
	.datab(!saved_grant_0),
	.datac(!\out_endofpacket~0_combout ),
	.datad(!nxt_in_ready2),
	.datae(!\use_reg~q ),
	.dataf(!nxt_in_ready1),
	.datag(!src0_valid1),
	.cin(gnd),
	.sharein(gnd),
	.combout(\use_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \use_reg~0 .extended_lut = "on";
defparam \use_reg~0 .lut_mask = 64'h0001FFF00101F0F0;
defparam \use_reg~0 .shared_arith = "off";

dffeas use_reg(
	.clk(outclk_wire_0),
	.d(\use_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\use_reg~q ),
	.prn(vcc));
defparam use_reg.is_wysiwyg = "true";
defparam use_reg.power_up = "low";

cyclonev_lcell_comb \address_reg~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready),
	.datac(!out_valid_reg),
	.datad(!cp_ready),
	.datae(!\use_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\address_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \address_reg~0 .extended_lut = "off";
defparam \address_reg~0 .lut_mask = 64'hFFFFD1DDFFFFD1DD;
defparam \address_reg~0 .shared_arith = "off";

dffeas \address_reg[1] (
	.clk(outclk_wire_0),
	.d(\Add1~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\address_reg[1]~q ),
	.prn(vcc));
defparam \address_reg[1] .is_wysiwyg = "true";
defparam \address_reg[1] .power_up = "low";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!src_payload),
	.datab(!src_payload1),
	.datac(!src_payload2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'h1010101010101010;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!src_payload),
	.datab(!src_payload1),
	.datac(!src_payload2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'h4040404040404040;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!count_0),
	.datab(!\use_reg~q ),
	.datac(!\Decoder0~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'hE2E2E2E2E2E2E2E2;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!count_1),
	.datab(!\use_reg~q ),
	.datac(!\Decoder0~0_combout ),
	.datad(!\Add0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h1DE21DE21DE21DE2;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \count~0 (
	.dataa(!saved_grant_0),
	.datab(!LessThan2),
	.datac(!Equal0),
	.datad(!Equal01),
	.datae(!Equal02),
	.dataf(!src0_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~0 .extended_lut = "off";
defparam \count~0 .lut_mask = 64'h0000000000000001;
defparam \count~0 .shared_arith = "off";

cyclonev_lcell_comb \count~1 (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready),
	.datac(!out_valid_reg),
	.datad(!cp_ready),
	.datae(!\use_reg~q ),
	.dataf(!\count~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~1 .extended_lut = "off";
defparam \count~1 .lut_mask = 64'h0000D1DDD1DDD1DD;
defparam \count~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\LessThan3~0_combout ),
	.datab(!\Decoder0~2_combout ),
	.datac(!\Decoder0~3_combout ),
	.datad(!int_output_sel_0),
	.datae(gnd),
	.dataf(!\Decoder0~1_combout ),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h00008000000000FF;
defparam \Add1~1 .shared_arith = "off";

dffeas \address_reg[2] (
	.clk(outclk_wire_0),
	.d(\Add1~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\address_reg[2]~q ),
	.prn(vcc));
defparam \address_reg[2] .is_wysiwyg = "true";
defparam \address_reg[2] .power_up = "low";

cyclonev_lcell_comb \Add1~5 (
	.dataa(!\LessThan3~0_combout ),
	.datab(!\Decoder0~2_combout ),
	.datac(!\Decoder0~3_combout ),
	.datad(!int_output_sel_1),
	.datae(gnd),
	.dataf(!\Decoder0~0_combout ),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FF7F000000FF;
defparam \Add1~5 .shared_arith = "off";

dffeas \address_reg[3] (
	.clk(outclk_wire_0),
	.d(\Add1~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\address_reg[3]~q ),
	.prn(vcc));
defparam \address_reg[3] .is_wysiwyg = "true";
defparam \address_reg[3] .power_up = "low";

cyclonev_lcell_comb \endofpacket_reg~0 (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_0),
	.datac(!\use_reg~q ),
	.datad(!\endofpacket_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\endofpacket_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \endofpacket_reg~0 .extended_lut = "off";
defparam \endofpacket_reg~0 .lut_mask = 64'h101F101F101F101F;
defparam \endofpacket_reg~0 .shared_arith = "off";

dffeas endofpacket_reg(
	.clk(outclk_wire_0),
	.d(\endofpacket_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\endofpacket_reg~q ),
	.prn(vcc));
defparam endofpacket_reg.is_wysiwyg = "true";
defparam endofpacket_reg.power_up = "low";

dffeas \address_reg[0] (
	.clk(outclk_wire_0),
	.d(\Add1~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\address_reg[0]~q ),
	.prn(vcc));
defparam \address_reg[0] .is_wysiwyg = "true";
defparam \address_reg[0] .power_up = "low";

endmodule

module Computer_System_altera_merlin_width_adapter_1 (
	h2f_BREADY_0,
	h2f_RREADY_0,
	outclk_wire_0,
	data_reg_0,
	data_reg_32,
	data_reg_64,
	mem_68_0,
	mem_122_0,
	mem_123_0,
	mem_124_0,
	mem_90_0,
	mem_91_0,
	ShiftRight0,
	source_addr_2,
	always10,
	mem_126_0,
	source_addr_3,
	always101,
	mem_31_0,
	LessThan15,
	r_sync_rst,
	p1_ready,
	read,
	always102)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	outclk_wire_0;
output 	data_reg_0;
output 	data_reg_32;
output 	data_reg_64;
input 	mem_68_0;
input 	mem_122_0;
input 	mem_123_0;
input 	mem_124_0;
input 	mem_90_0;
input 	mem_91_0;
output 	ShiftRight0;
input 	source_addr_2;
output 	always10;
input 	mem_126_0;
input 	source_addr_3;
output 	always101;
input 	mem_31_0;
output 	LessThan15;
input 	r_sync_rst;
output 	p1_ready;
input 	read;
output 	always102;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_reg~0_combout ;
wire \data_reg~1_combout ;
wire \data_reg~2_combout ;


dffeas \data_reg[0] (
	.clk(outclk_wire_0),
	.d(\data_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always102),
	.sload(gnd),
	.ena(read),
	.q(data_reg_0),
	.prn(vcc));
defparam \data_reg[0] .is_wysiwyg = "true";
defparam \data_reg[0] .power_up = "low";

dffeas \data_reg[32] (
	.clk(outclk_wire_0),
	.d(\data_reg~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always102),
	.sload(gnd),
	.ena(read),
	.q(data_reg_32),
	.prn(vcc));
defparam \data_reg[32] .is_wysiwyg = "true";
defparam \data_reg[32] .power_up = "low";

dffeas \data_reg[64] (
	.clk(outclk_wire_0),
	.d(\data_reg~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always102),
	.sload(gnd),
	.ena(read),
	.q(data_reg_64),
	.prn(vcc));
defparam \data_reg[64] .is_wysiwyg = "true";
defparam \data_reg[64] .power_up = "low";

cyclonev_lcell_comb \ShiftRight0~0 (
	.dataa(!mem_122_0),
	.datab(!mem_123_0),
	.datac(!mem_124_0),
	.datad(!mem_90_0),
	.datae(!mem_91_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftRight0),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftRight0~0 .extended_lut = "off";
defparam \ShiftRight0~0 .lut_mask = 64'h0804020108040201;
defparam \ShiftRight0~0 .shared_arith = "off";

cyclonev_lcell_comb \always10~0 (
	.dataa(!source_addr_2),
	.datab(!mem_122_0),
	.datac(!mem_123_0),
	.datad(!mem_124_0),
	.datae(!mem_90_0),
	.dataf(!mem_91_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always10),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~0 .extended_lut = "off";
defparam \always10~0 .lut_mask = 64'hE0C0F830FE0CFF83;
defparam \always10~0 .shared_arith = "off";

cyclonev_lcell_comb \always10~1 (
	.dataa(!mem_126_0),
	.datab(!source_addr_2),
	.datac(!source_addr_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always101),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~1 .extended_lut = "off";
defparam \always10~1 .lut_mask = 64'h2A2A2A2A2A2A2A2A;
defparam \always10~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan15~0 (
	.dataa(!mem_122_0),
	.datab(!mem_123_0),
	.datac(!mem_124_0),
	.datad(!mem_90_0),
	.datae(!mem_91_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan15),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan15~0 .extended_lut = "off";
defparam \LessThan15~0 .lut_mask = 64'h80C0E0F080C0E0F0;
defparam \LessThan15~0 .shared_arith = "off";

cyclonev_lcell_comb \p1_ready~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!h2f_RREADY_0),
	.datac(!mem_68_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(p1_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_ready~0 .extended_lut = "off";
defparam \p1_ready~0 .lut_mask = 64'h3535353535353535;
defparam \p1_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \always10~2 (
	.dataa(!ShiftRight0),
	.datab(!always10),
	.datac(!always101),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always102),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~2 .extended_lut = "off";
defparam \always10~2 .lut_mask = 64'hF2F2F2F2F2F2F2F2;
defparam \always10~2 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~0 (
	.dataa(!source_addr_2),
	.datab(!source_addr_3),
	.datac(!mem_31_0),
	.datad(!data_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~0 .extended_lut = "off";
defparam \data_reg~0 .lut_mask = 64'h01FF01FF01FF01FF;
defparam \data_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~1 (
	.dataa(!source_addr_2),
	.datab(!source_addr_3),
	.datac(!mem_31_0),
	.datad(!data_reg_32),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~1 .extended_lut = "off";
defparam \data_reg~1 .lut_mask = 64'h02FF02FF02FF02FF;
defparam \data_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~2 (
	.dataa(!source_addr_2),
	.datab(!source_addr_3),
	.datac(!mem_31_0),
	.datad(!data_reg_64),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~2 .extended_lut = "off";
defparam \data_reg~2 .lut_mask = 64'h04FF04FF04FF04FF;
defparam \data_reg~2 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_width_adapter_2 (
	h2f_WLAST_0,
	h2f_ARADDR_1,
	h2f_ARADDR_3,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWADDR_1,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WDATA_0,
	h2f_WDATA_1,
	h2f_WDATA_2,
	h2f_WDATA_3,
	h2f_WDATA_4,
	h2f_WDATA_5,
	h2f_WDATA_6,
	h2f_WDATA_7,
	h2f_WDATA_8,
	h2f_WDATA_9,
	h2f_WDATA_10,
	h2f_WDATA_11,
	h2f_WDATA_12,
	h2f_WDATA_13,
	h2f_WDATA_14,
	h2f_WDATA_15,
	h2f_WDATA_16,
	h2f_WDATA_17,
	h2f_WDATA_18,
	h2f_WDATA_19,
	h2f_WDATA_20,
	h2f_WDATA_21,
	h2f_WDATA_22,
	h2f_WDATA_23,
	h2f_WDATA_24,
	h2f_WDATA_25,
	h2f_WDATA_26,
	h2f_WDATA_27,
	h2f_WDATA_28,
	h2f_WDATA_29,
	h2f_WDATA_30,
	h2f_WDATA_31,
	h2f_WDATA_32,
	h2f_WDATA_33,
	h2f_WDATA_34,
	h2f_WDATA_35,
	h2f_WDATA_36,
	h2f_WDATA_37,
	h2f_WDATA_38,
	h2f_WDATA_39,
	h2f_WDATA_40,
	h2f_WDATA_41,
	h2f_WDATA_42,
	h2f_WDATA_43,
	h2f_WDATA_44,
	h2f_WDATA_45,
	h2f_WDATA_46,
	h2f_WDATA_47,
	h2f_WDATA_48,
	h2f_WDATA_49,
	h2f_WDATA_50,
	h2f_WDATA_51,
	h2f_WDATA_52,
	h2f_WDATA_53,
	h2f_WDATA_54,
	h2f_WDATA_55,
	h2f_WDATA_56,
	h2f_WDATA_57,
	h2f_WDATA_58,
	h2f_WDATA_59,
	h2f_WDATA_60,
	h2f_WDATA_61,
	h2f_WDATA_62,
	h2f_WDATA_63,
	h2f_WDATA_64,
	h2f_WDATA_65,
	h2f_WDATA_66,
	h2f_WDATA_67,
	h2f_WDATA_68,
	h2f_WDATA_69,
	h2f_WDATA_70,
	h2f_WDATA_71,
	h2f_WDATA_72,
	h2f_WDATA_73,
	h2f_WDATA_74,
	h2f_WDATA_75,
	h2f_WDATA_76,
	h2f_WDATA_77,
	h2f_WDATA_78,
	h2f_WDATA_79,
	h2f_WDATA_80,
	h2f_WDATA_81,
	h2f_WDATA_82,
	h2f_WDATA_83,
	h2f_WDATA_84,
	h2f_WDATA_85,
	h2f_WDATA_86,
	h2f_WDATA_87,
	h2f_WDATA_88,
	h2f_WDATA_89,
	h2f_WDATA_90,
	h2f_WDATA_91,
	h2f_WDATA_92,
	h2f_WDATA_93,
	h2f_WDATA_94,
	h2f_WDATA_95,
	h2f_WDATA_96,
	h2f_WDATA_97,
	h2f_WDATA_98,
	h2f_WDATA_99,
	h2f_WDATA_100,
	h2f_WDATA_101,
	h2f_WDATA_102,
	h2f_WDATA_103,
	h2f_WDATA_104,
	h2f_WDATA_105,
	h2f_WDATA_106,
	h2f_WDATA_107,
	h2f_WDATA_108,
	h2f_WDATA_109,
	h2f_WDATA_110,
	h2f_WDATA_111,
	h2f_WDATA_112,
	h2f_WDATA_113,
	h2f_WDATA_114,
	h2f_WDATA_115,
	h2f_WDATA_116,
	h2f_WDATA_117,
	h2f_WDATA_118,
	h2f_WDATA_119,
	h2f_WDATA_120,
	h2f_WDATA_121,
	h2f_WDATA_122,
	h2f_WDATA_123,
	h2f_WDATA_124,
	h2f_WDATA_125,
	h2f_WDATA_126,
	h2f_WDATA_127,
	outclk_wire_0,
	Mux4,
	Mux5,
	Mux6,
	Mux7,
	Mux8,
	Mux9,
	Mux10,
	Mux11,
	Mux12,
	Mux13,
	Mux14,
	Mux15,
	Mux16,
	Mux17,
	Mux18,
	Mux19,
	Mux20,
	Mux21,
	Mux22,
	Mux23,
	Mux24,
	Mux25,
	Mux26,
	Mux27,
	Mux28,
	Mux29,
	Mux30,
	Mux31,
	Mux32,
	Mux33,
	Mux34,
	Mux35,
	src_data_185,
	saved_grant_1,
	saved_grant_0,
	src_data_198,
	src_data_199,
	src_data_200,
	in_ready,
	nxt_in_ready,
	nxt_in_ready1,
	sop_enable,
	r_sync_rst,
	WideOr1,
	in_endofpacket,
	use_reg1,
	out_data_91,
	out_data_90,
	address_burst_1,
	out_data_37,
	src_data_144,
	out_data_36,
	src_data_130,
	src_data_134,
	src_data_138,
	src_data_142,
	src_data_146,
	int_output_sel_0,
	out_data_3,
	Mux1,
	src_data_128,
	src_data_132,
	src_data_136,
	src_data_140,
	Mux3,
	src_data_129,
	src_data_133,
	src_data_137,
	src_data_141,
	Mux2,
	src_data_131,
	src_data_135,
	src_data_139,
	src_data_143,
	Mux0,
	out_endofpacket,
	src_data_184,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	out_data_74,
	src_data_187,
	src_data_186,
	write_cp_data_188,
	src_payload4,
	src_data_188,
	out_data_79,
	out_data_76,
	write_cp_data_187,
	src_payload5,
	out_data_77,
	out_data_78,
	out_data_80,
	out_data_75,
	out_data_7,
	out_data_6,
	out_data_4,
	out_data_5,
	address_reg_4,
	src_payload6,
	address_reg_5,
	src_payload7,
	address_reg_6,
	src_payload8,
	address_reg_7,
	src_payload9,
	src_data_152,
	out_data_44,
	src_payload10,
	src_payload11,
	out_data_45,
	int_output_sel_1)/* synthesis synthesis_greybox=0 */;
input 	h2f_WLAST_0;
input 	h2f_ARADDR_1;
input 	h2f_ARADDR_3;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWADDR_1;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WDATA_0;
input 	h2f_WDATA_1;
input 	h2f_WDATA_2;
input 	h2f_WDATA_3;
input 	h2f_WDATA_4;
input 	h2f_WDATA_5;
input 	h2f_WDATA_6;
input 	h2f_WDATA_7;
input 	h2f_WDATA_8;
input 	h2f_WDATA_9;
input 	h2f_WDATA_10;
input 	h2f_WDATA_11;
input 	h2f_WDATA_12;
input 	h2f_WDATA_13;
input 	h2f_WDATA_14;
input 	h2f_WDATA_15;
input 	h2f_WDATA_16;
input 	h2f_WDATA_17;
input 	h2f_WDATA_18;
input 	h2f_WDATA_19;
input 	h2f_WDATA_20;
input 	h2f_WDATA_21;
input 	h2f_WDATA_22;
input 	h2f_WDATA_23;
input 	h2f_WDATA_24;
input 	h2f_WDATA_25;
input 	h2f_WDATA_26;
input 	h2f_WDATA_27;
input 	h2f_WDATA_28;
input 	h2f_WDATA_29;
input 	h2f_WDATA_30;
input 	h2f_WDATA_31;
input 	h2f_WDATA_32;
input 	h2f_WDATA_33;
input 	h2f_WDATA_34;
input 	h2f_WDATA_35;
input 	h2f_WDATA_36;
input 	h2f_WDATA_37;
input 	h2f_WDATA_38;
input 	h2f_WDATA_39;
input 	h2f_WDATA_40;
input 	h2f_WDATA_41;
input 	h2f_WDATA_42;
input 	h2f_WDATA_43;
input 	h2f_WDATA_44;
input 	h2f_WDATA_45;
input 	h2f_WDATA_46;
input 	h2f_WDATA_47;
input 	h2f_WDATA_48;
input 	h2f_WDATA_49;
input 	h2f_WDATA_50;
input 	h2f_WDATA_51;
input 	h2f_WDATA_52;
input 	h2f_WDATA_53;
input 	h2f_WDATA_54;
input 	h2f_WDATA_55;
input 	h2f_WDATA_56;
input 	h2f_WDATA_57;
input 	h2f_WDATA_58;
input 	h2f_WDATA_59;
input 	h2f_WDATA_60;
input 	h2f_WDATA_61;
input 	h2f_WDATA_62;
input 	h2f_WDATA_63;
input 	h2f_WDATA_64;
input 	h2f_WDATA_65;
input 	h2f_WDATA_66;
input 	h2f_WDATA_67;
input 	h2f_WDATA_68;
input 	h2f_WDATA_69;
input 	h2f_WDATA_70;
input 	h2f_WDATA_71;
input 	h2f_WDATA_72;
input 	h2f_WDATA_73;
input 	h2f_WDATA_74;
input 	h2f_WDATA_75;
input 	h2f_WDATA_76;
input 	h2f_WDATA_77;
input 	h2f_WDATA_78;
input 	h2f_WDATA_79;
input 	h2f_WDATA_80;
input 	h2f_WDATA_81;
input 	h2f_WDATA_82;
input 	h2f_WDATA_83;
input 	h2f_WDATA_84;
input 	h2f_WDATA_85;
input 	h2f_WDATA_86;
input 	h2f_WDATA_87;
input 	h2f_WDATA_88;
input 	h2f_WDATA_89;
input 	h2f_WDATA_90;
input 	h2f_WDATA_91;
input 	h2f_WDATA_92;
input 	h2f_WDATA_93;
input 	h2f_WDATA_94;
input 	h2f_WDATA_95;
input 	h2f_WDATA_96;
input 	h2f_WDATA_97;
input 	h2f_WDATA_98;
input 	h2f_WDATA_99;
input 	h2f_WDATA_100;
input 	h2f_WDATA_101;
input 	h2f_WDATA_102;
input 	h2f_WDATA_103;
input 	h2f_WDATA_104;
input 	h2f_WDATA_105;
input 	h2f_WDATA_106;
input 	h2f_WDATA_107;
input 	h2f_WDATA_108;
input 	h2f_WDATA_109;
input 	h2f_WDATA_110;
input 	h2f_WDATA_111;
input 	h2f_WDATA_112;
input 	h2f_WDATA_113;
input 	h2f_WDATA_114;
input 	h2f_WDATA_115;
input 	h2f_WDATA_116;
input 	h2f_WDATA_117;
input 	h2f_WDATA_118;
input 	h2f_WDATA_119;
input 	h2f_WDATA_120;
input 	h2f_WDATA_121;
input 	h2f_WDATA_122;
input 	h2f_WDATA_123;
input 	h2f_WDATA_124;
input 	h2f_WDATA_125;
input 	h2f_WDATA_126;
input 	h2f_WDATA_127;
input 	outclk_wire_0;
output 	Mux4;
output 	Mux5;
output 	Mux6;
output 	Mux7;
output 	Mux8;
output 	Mux9;
output 	Mux10;
output 	Mux11;
output 	Mux12;
output 	Mux13;
output 	Mux14;
output 	Mux15;
output 	Mux16;
output 	Mux17;
output 	Mux18;
output 	Mux19;
output 	Mux20;
output 	Mux21;
output 	Mux22;
output 	Mux23;
output 	Mux24;
output 	Mux25;
output 	Mux26;
output 	Mux27;
output 	Mux28;
output 	Mux29;
output 	Mux30;
output 	Mux31;
output 	Mux32;
output 	Mux33;
output 	Mux34;
output 	Mux35;
input 	src_data_185;
input 	saved_grant_1;
input 	saved_grant_0;
input 	src_data_198;
input 	src_data_199;
input 	src_data_200;
output 	in_ready;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	sop_enable;
input 	r_sync_rst;
input 	WideOr1;
input 	in_endofpacket;
output 	use_reg1;
output 	out_data_91;
output 	out_data_90;
input 	address_burst_1;
output 	out_data_37;
input 	src_data_144;
output 	out_data_36;
input 	src_data_130;
input 	src_data_134;
input 	src_data_138;
input 	src_data_142;
input 	src_data_146;
output 	int_output_sel_0;
input 	out_data_3;
output 	Mux1;
input 	src_data_128;
input 	src_data_132;
input 	src_data_136;
input 	src_data_140;
output 	Mux3;
input 	src_data_129;
input 	src_data_133;
input 	src_data_137;
input 	src_data_141;
output 	Mux2;
input 	src_data_131;
input 	src_data_135;
input 	src_data_139;
input 	src_data_143;
output 	Mux0;
output 	out_endofpacket;
input 	src_data_184;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
output 	out_data_74;
input 	src_data_187;
input 	src_data_186;
input 	write_cp_data_188;
input 	src_payload4;
input 	src_data_188;
output 	out_data_79;
output 	out_data_76;
input 	write_cp_data_187;
input 	src_payload5;
output 	out_data_77;
output 	out_data_78;
output 	out_data_80;
output 	out_data_75;
input 	out_data_7;
input 	out_data_6;
input 	out_data_4;
input 	out_data_5;
output 	address_reg_4;
input 	src_payload6;
output 	address_reg_5;
input 	src_payload7;
output 	address_reg_6;
input 	src_payload8;
output 	address_reg_7;
input 	src_payload9;
input 	src_data_152;
output 	out_data_44;
input 	src_payload10;
input 	src_payload11;
output 	out_data_45;
output 	int_output_sel_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Decoder0~0_combout ;
wire \in_ready~1_combout ;
wire \count~0_combout ;
wire \count[0]~q ;
wire \Decoder0~1_combout ;
wire \Add0~0_combout ;
wire \Add0~1_combout ;
wire \count[1]~q ;
wire \out_endofpacket~0_combout ;
wire \use_reg~0_combout ;
wire \Decoder0~3_combout ;
wire \Decoder0~4_combout ;
wire \Decoder0~2_combout ;
wire \Decoder0~5_combout ;
wire \LessThan3~0_combout ;
wire \Decoder0~6_combout ;
wire \Add1~6 ;
wire \Add1~1_sumout ;
wire \address_reg~0_combout ;
wire \address_reg[1]~q ;
wire \out_data[37]~2_combout ;
wire \Add1~5_sumout ;
wire \address_reg[0]~q ;
wire \Add1~2 ;
wire \Add1~9_sumout ;
wire \address_reg[2]~q ;
wire \endofpacket_reg~q ;
wire \LessThan2~0_combout ;
wire \out_endofpacket~1_combout ;
wire \ShiftLeft0~6_combout ;
wire \byte_cnt_reg~0_combout ;
wire \byte_cnt_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \int_byte_cnt_factor[0]~0_combout ;
wire \ShiftLeft0~2_combout ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~7_combout ;
wire \ShiftLeft0~1_combout ;
wire \out_data[78]~12_combout ;
wire \out_data[78]~13_combout ;
wire \out_data[78]~20_combout ;
wire \out_data[77]~8_combout ;
wire \out_data[77]~9_combout ;
wire \out_data[77]~10_combout ;
wire \out_data[77]~19_combout ;
wire \ShiftLeft0~4_combout ;
wire \ShiftLeft0~5_combout ;
wire \ShiftLeft0~8_combout ;
wire \Add2~26_cout ;
wire \Add2~21_sumout ;
wire \byte_cnt_reg[3]~q ;
wire \Add2~22 ;
wire \Add2~5_sumout ;
wire \byte_cnt_reg[4]~q ;
wire \Add2~6 ;
wire \Add2~9_sumout ;
wire \byte_cnt_reg[5]~q ;
wire \Add2~10 ;
wire \Add2~13_sumout ;
wire \byte_cnt_reg[6]~q ;
wire \Add2~14 ;
wire \Add2~1_sumout ;
wire \byte_cnt_reg[7]~q ;
wire \Add2~2 ;
wire \Add2~17_sumout ;
wire \byte_cnt_reg[8]~q ;
wire \Add1~10 ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \Add1~22 ;
wire \Add1~25_sumout ;
wire \Add1~26 ;
wire \Add1~29_sumout ;
wire \Add1~30 ;
wire \Add1~33_sumout ;
wire \address_reg[8]~q ;
wire \Add1~34 ;
wire \Add1~37_sumout ;
wire \address_reg[9]~q ;
wire \int_output_sel[1]~1_combout ;
wire \Add1~13_sumout ;
wire \address_reg[3]~q ;


cyclonev_lcell_comb \Mux4~0 (
	.dataa(!h2f_WDATA_127),
	.datab(!h2f_WDATA_63),
	.datac(!h2f_WDATA_95),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_31),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~0 .extended_lut = "on";
defparam \Mux4~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux4~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux5~0 (
	.dataa(!h2f_WDATA_126),
	.datab(!h2f_WDATA_62),
	.datac(!h2f_WDATA_94),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_30),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux5),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~0 .extended_lut = "on";
defparam \Mux5~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux5~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux6~0 (
	.dataa(!h2f_WDATA_125),
	.datab(!h2f_WDATA_61),
	.datac(!h2f_WDATA_93),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_29),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux6),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~0 .extended_lut = "on";
defparam \Mux6~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux6~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux7~0 (
	.dataa(!h2f_WDATA_124),
	.datab(!h2f_WDATA_60),
	.datac(!h2f_WDATA_92),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_28),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux7),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~0 .extended_lut = "on";
defparam \Mux7~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux7~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~0 (
	.dataa(!h2f_WDATA_123),
	.datab(!h2f_WDATA_59),
	.datac(!h2f_WDATA_91),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_27),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux8),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~0 .extended_lut = "on";
defparam \Mux8~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux8~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux9~0 (
	.dataa(!h2f_WDATA_122),
	.datab(!h2f_WDATA_58),
	.datac(!h2f_WDATA_90),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_26),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux9),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~0 .extended_lut = "on";
defparam \Mux9~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux9~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux10~0 (
	.dataa(!h2f_WDATA_121),
	.datab(!h2f_WDATA_57),
	.datac(!h2f_WDATA_89),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_25),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux10),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~0 .extended_lut = "on";
defparam \Mux10~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux10~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux11~0 (
	.dataa(!h2f_WDATA_120),
	.datab(!h2f_WDATA_56),
	.datac(!h2f_WDATA_88),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_24),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~0 .extended_lut = "on";
defparam \Mux11~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux11~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux12~0 (
	.dataa(!h2f_WDATA_119),
	.datab(!h2f_WDATA_55),
	.datac(!h2f_WDATA_87),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_23),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux12),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux12~0 .extended_lut = "on";
defparam \Mux12~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux12~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux13~0 (
	.dataa(!h2f_WDATA_118),
	.datab(!h2f_WDATA_54),
	.datac(!h2f_WDATA_86),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_22),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux13),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~0 .extended_lut = "on";
defparam \Mux13~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux13~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux14~0 (
	.dataa(!h2f_WDATA_117),
	.datab(!h2f_WDATA_53),
	.datac(!h2f_WDATA_85),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_21),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux14),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~0 .extended_lut = "on";
defparam \Mux14~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux14~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux15~0 (
	.dataa(!h2f_WDATA_116),
	.datab(!h2f_WDATA_52),
	.datac(!h2f_WDATA_84),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_20),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux15),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux15~0 .extended_lut = "on";
defparam \Mux15~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux15~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux16~0 (
	.dataa(!h2f_WDATA_115),
	.datab(!h2f_WDATA_51),
	.datac(!h2f_WDATA_83),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_19),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux16),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~0 .extended_lut = "on";
defparam \Mux16~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux16~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux17~0 (
	.dataa(!h2f_WDATA_114),
	.datab(!h2f_WDATA_50),
	.datac(!h2f_WDATA_82),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_18),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux17),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux17~0 .extended_lut = "on";
defparam \Mux17~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux17~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux18~0 (
	.dataa(!h2f_WDATA_113),
	.datab(!h2f_WDATA_49),
	.datac(!h2f_WDATA_81),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_17),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux18),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux18~0 .extended_lut = "on";
defparam \Mux18~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux18~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux19~0 (
	.dataa(!h2f_WDATA_112),
	.datab(!h2f_WDATA_48),
	.datac(!h2f_WDATA_80),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_16),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux19),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux19~0 .extended_lut = "on";
defparam \Mux19~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux19~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux20~0 (
	.dataa(!h2f_WDATA_111),
	.datab(!h2f_WDATA_47),
	.datac(!h2f_WDATA_79),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_15),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux20),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux20~0 .extended_lut = "on";
defparam \Mux20~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux20~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux21~0 (
	.dataa(!h2f_WDATA_110),
	.datab(!h2f_WDATA_46),
	.datac(!h2f_WDATA_78),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_14),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux21),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux21~0 .extended_lut = "on";
defparam \Mux21~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux21~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux22~0 (
	.dataa(!h2f_WDATA_109),
	.datab(!h2f_WDATA_45),
	.datac(!h2f_WDATA_77),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_13),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux22),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~0 .extended_lut = "on";
defparam \Mux22~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux22~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux23~0 (
	.dataa(!h2f_WDATA_108),
	.datab(!h2f_WDATA_44),
	.datac(!h2f_WDATA_76),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_12),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux23),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux23~0 .extended_lut = "on";
defparam \Mux23~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux23~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~0 (
	.dataa(!h2f_WDATA_107),
	.datab(!h2f_WDATA_43),
	.datac(!h2f_WDATA_75),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_11),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux24),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~0 .extended_lut = "on";
defparam \Mux24~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux24~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux25~0 (
	.dataa(!h2f_WDATA_106),
	.datab(!h2f_WDATA_42),
	.datac(!h2f_WDATA_74),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_10),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux25),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~0 .extended_lut = "on";
defparam \Mux25~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux25~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux26~0 (
	.dataa(!h2f_WDATA_105),
	.datab(!h2f_WDATA_41),
	.datac(!h2f_WDATA_73),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_9),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux26),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~0 .extended_lut = "on";
defparam \Mux26~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux26~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux27~0 (
	.dataa(!h2f_WDATA_104),
	.datab(!h2f_WDATA_40),
	.datac(!h2f_WDATA_72),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_8),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux27),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~0 .extended_lut = "on";
defparam \Mux27~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux27~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux28~0 (
	.dataa(!h2f_WDATA_103),
	.datab(!h2f_WDATA_39),
	.datac(!h2f_WDATA_71),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_7),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux28),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux28~0 .extended_lut = "on";
defparam \Mux28~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux28~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux29~0 (
	.dataa(!h2f_WDATA_102),
	.datab(!h2f_WDATA_38),
	.datac(!h2f_WDATA_70),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_6),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux29),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux29~0 .extended_lut = "on";
defparam \Mux29~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux29~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux30~0 (
	.dataa(!h2f_WDATA_101),
	.datab(!h2f_WDATA_37),
	.datac(!h2f_WDATA_69),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_5),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux30),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux30~0 .extended_lut = "on";
defparam \Mux30~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux30~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux31~0 (
	.dataa(!h2f_WDATA_100),
	.datab(!h2f_WDATA_36),
	.datac(!h2f_WDATA_68),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_4),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux31),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux31~0 .extended_lut = "on";
defparam \Mux31~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux31~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~0 (
	.dataa(!h2f_WDATA_99),
	.datab(!h2f_WDATA_35),
	.datac(!h2f_WDATA_67),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_3),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux32),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~0 .extended_lut = "on";
defparam \Mux32~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux32~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux33~0 (
	.dataa(!h2f_WDATA_98),
	.datab(!h2f_WDATA_34),
	.datac(!h2f_WDATA_66),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_2),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux33),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux33~0 .extended_lut = "on";
defparam \Mux33~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux33~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux34~0 (
	.dataa(!h2f_WDATA_97),
	.datab(!h2f_WDATA_33),
	.datac(!h2f_WDATA_65),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux34),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux34~0 .extended_lut = "on";
defparam \Mux34~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux34~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux35~0 (
	.dataa(!h2f_WDATA_96),
	.datab(!h2f_WDATA_32),
	.datac(!h2f_WDATA_64),
	.datad(!saved_grant_0),
	.datae(!int_output_sel_1),
	.dataf(!int_output_sel_0),
	.datag(!h2f_WDATA_0),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux35),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux35~0 .extended_lut = "on";
defparam \Mux35~0 .lut_mask = 64'h000F000F00330055;
defparam \Mux35~0 .shared_arith = "off";

cyclonev_lcell_comb \in_ready~0 (
	.dataa(!saved_grant_1),
	.datab(!\out_endofpacket~0_combout ),
	.datac(!src_data_198),
	.datad(!src_data_199),
	.datae(!src_data_200),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_ready~0 .extended_lut = "off";
defparam \in_ready~0 .lut_mask = 64'h0008888800088888;
defparam \in_ready~0 .shared_arith = "off";

dffeas use_reg(
	.clk(outclk_wire_0),
	.d(\use_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(use_reg1),
	.prn(vcc));
defparam use_reg.is_wysiwyg = "true";
defparam use_reg.power_up = "low";

cyclonev_lcell_comb \out_data[91]~0 (
	.dataa(!src_data_199),
	.datab(!src_data_200),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_91),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[91]~0 .extended_lut = "off";
defparam \out_data[91]~0 .lut_mask = 64'h7777777777777777;
defparam \out_data[91]~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[90]~1 (
	.dataa(!src_data_198),
	.datab(!src_data_199),
	.datac(!src_data_200),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_90),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[90]~1 .extended_lut = "off";
defparam \out_data[90]~1 .lut_mask = 64'h4040404040404040;
defparam \out_data[90]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[37]~3 (
	.dataa(!src_data_198),
	.datab(!src_data_199),
	.datac(!src_data_200),
	.datad(!use_reg1),
	.datae(!\address_reg[1]~q ),
	.dataf(!\out_data[37]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_37),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[37]~3 .extended_lut = "off";
defparam \out_data[37]~3 .lut_mask = 64'h000000FFE000E0FF;
defparam \out_data[37]~3 .shared_arith = "off";

cyclonev_lcell_comb \out_data[36]~4 (
	.dataa(!src_data_198),
	.datab(!src_data_199),
	.datac(!src_data_200),
	.datad(!use_reg1),
	.datae(!\address_reg[0]~q ),
	.dataf(!src_data_144),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_36),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[36]~4 .extended_lut = "off";
defparam \out_data[36]~4 .lut_mask = 64'h000000FFE000E0FF;
defparam \out_data[36]~4 .shared_arith = "off";

cyclonev_lcell_comb \int_output_sel[0]~0 (
	.dataa(!src_data_198),
	.datab(!src_data_199),
	.datac(!src_data_200),
	.datad(!use_reg1),
	.datae(!\address_reg[2]~q ),
	.dataf(!src_data_146),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(int_output_sel_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_output_sel[0]~0 .extended_lut = "off";
defparam \int_output_sel[0]~0 .lut_mask = 64'h000000FFE000E0FF;
defparam \int_output_sel[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux1~0 (
	.dataa(!src_data_130),
	.datab(!src_data_134),
	.datac(!src_data_138),
	.datad(!src_data_142),
	.datae(!int_output_sel_0),
	.dataf(!int_output_sel_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~0 .extended_lut = "off";
defparam \Mux1~0 .lut_mask = 64'hAAAACCCCF0F0FF00;
defparam \Mux1~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~0 (
	.dataa(!src_data_128),
	.datab(!src_data_132),
	.datac(!src_data_136),
	.datad(!src_data_140),
	.datae(!int_output_sel_0),
	.dataf(!int_output_sel_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'hAAAACCCCF0F0FF00;
defparam \Mux3~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~0 (
	.dataa(!src_data_129),
	.datab(!src_data_133),
	.datac(!src_data_137),
	.datad(!src_data_141),
	.datae(!int_output_sel_0),
	.dataf(!int_output_sel_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~0 .extended_lut = "off";
defparam \Mux2~0 .lut_mask = 64'hAAAACCCCF0F0FF00;
defparam \Mux2~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!src_data_131),
	.datab(!src_data_135),
	.datac(!src_data_139),
	.datad(!src_data_143),
	.datae(!int_output_sel_0),
	.dataf(!int_output_sel_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'hAAAACCCCF0F0FF00;
defparam \Mux0~0 .shared_arith = "off";

cyclonev_lcell_comb \out_endofpacket~2 (
	.dataa(!\out_endofpacket~0_combout ),
	.datab(!use_reg1),
	.datac(!\endofpacket_reg~q ),
	.datad(!\out_endofpacket~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_endofpacket),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_endofpacket~2 .extended_lut = "off";
defparam \out_endofpacket~2 .lut_mask = 64'hEF01EF01EF01EF01;
defparam \out_endofpacket~2 .shared_arith = "off";

cyclonev_lcell_comb \out_data[74]~5 (
	.dataa(gnd),
	.datab(!src_data_200),
	.datac(!use_reg1),
	.datad(!\byte_cnt_reg[2]~q ),
	.datae(!\ShiftLeft0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_74),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[74]~5 .extended_lut = "off";
defparam \out_data[74]~5 .lut_mask = 64'h000FC0CF000FC0CF;
defparam \out_data[74]~5 .shared_arith = "off";

cyclonev_lcell_comb \out_data[79]~6 (
	.dataa(!src_data_200),
	.datab(!\Decoder0~0_combout ),
	.datac(!use_reg1),
	.datad(!\byte_cnt_reg[7]~q ),
	.datae(!\ShiftLeft0~3_combout ),
	.dataf(!src_data_188),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[79]~6 .extended_lut = "off";
defparam \out_data[79]~6 .lut_mask = 64'h303F707F000F505F;
defparam \out_data[79]~6 .shared_arith = "off";

cyclonev_lcell_comb \out_data[76]~7 (
	.dataa(!src_data_200),
	.datab(!use_reg1),
	.datac(!\byte_cnt_reg[4]~q ),
	.datad(!\ShiftLeft0~4_combout ),
	.datae(!\ShiftLeft0~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_76),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[76]~7 .extended_lut = "off";
defparam \out_data[76]~7 .lut_mask = 64'h03CF8BCF03CF8BCF;
defparam \out_data[76]~7 .shared_arith = "off";

cyclonev_lcell_comb \out_data[77]~11 (
	.dataa(!src_data_200),
	.datab(!use_reg1),
	.datac(!\byte_cnt_reg[5]~q ),
	.datad(!\out_data[77]~8_combout ),
	.datae(!\out_data[77]~9_combout ),
	.dataf(!\out_data[77]~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_77),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[77]~11 .extended_lut = "off";
defparam \out_data[77]~11 .lut_mask = 64'h03CF8BCF8BCF8BCF;
defparam \out_data[77]~11 .shared_arith = "off";

cyclonev_lcell_comb \out_data[78]~14 (
	.dataa(!src_data_200),
	.datab(!use_reg1),
	.datac(!\ShiftLeft0~6_combout ),
	.datad(!\byte_cnt_reg[6]~q ),
	.datae(!\out_data[78]~12_combout ),
	.dataf(!\out_data[78]~13_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_78),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[78]~14 .extended_lut = "off";
defparam \out_data[78]~14 .lut_mask = 64'h04378CBF8CBF8CBF;
defparam \out_data[78]~14 .shared_arith = "off";

cyclonev_lcell_comb \out_data[80]~15 (
	.dataa(!src_data_200),
	.datab(!use_reg1),
	.datac(!\ShiftLeft0~5_combout ),
	.datad(!\byte_cnt_reg[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_80),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[80]~15 .extended_lut = "off";
defparam \out_data[80]~15 .lut_mask = 64'h0437043704370437;
defparam \out_data[80]~15 .shared_arith = "off";

cyclonev_lcell_comb \out_data[75]~16 (
	.dataa(!src_data_200),
	.datab(!use_reg1),
	.datac(!\ShiftLeft0~3_combout ),
	.datad(!\byte_cnt_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_75),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[75]~16 .extended_lut = "off";
defparam \out_data[75]~16 .lut_mask = 64'h083B083B083B083B;
defparam \out_data[75]~16 .shared_arith = "off";

dffeas \address_reg[4] (
	.clk(outclk_wire_0),
	.d(\Add1~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(address_reg_4),
	.prn(vcc));
defparam \address_reg[4] .is_wysiwyg = "true";
defparam \address_reg[4] .power_up = "low";

dffeas \address_reg[5] (
	.clk(outclk_wire_0),
	.d(\Add1~21_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(address_reg_5),
	.prn(vcc));
defparam \address_reg[5] .is_wysiwyg = "true";
defparam \address_reg[5] .power_up = "low";

dffeas \address_reg[6] (
	.clk(outclk_wire_0),
	.d(\Add1~25_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(address_reg_6),
	.prn(vcc));
defparam \address_reg[6] .is_wysiwyg = "true";
defparam \address_reg[6] .power_up = "low";

dffeas \address_reg[7] (
	.clk(outclk_wire_0),
	.d(\Add1~29_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(address_reg_7),
	.prn(vcc));
defparam \address_reg[7] .is_wysiwyg = "true";
defparam \address_reg[7] .power_up = "low";

cyclonev_lcell_comb \out_data[44]~17 (
	.dataa(!use_reg1),
	.datab(!\address_reg[8]~q ),
	.datac(!src_data_152),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[44]~17 .extended_lut = "off";
defparam \out_data[44]~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \out_data[44]~17 .shared_arith = "off";

cyclonev_lcell_comb \out_data[45]~18 (
	.dataa(!use_reg1),
	.datab(!\address_reg[9]~q ),
	.datac(!src_payload10),
	.datad(!src_payload11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[45]~18 .extended_lut = "off";
defparam \out_data[45]~18 .lut_mask = 64'h1BBB1BBB1BBB1BBB;
defparam \out_data[45]~18 .shared_arith = "off";

cyclonev_lcell_comb \int_output_sel[1]~2 (
	.dataa(!\int_output_sel[1]~1_combout ),
	.datab(!\address_reg[3]~q ),
	.datac(!use_reg1),
	.datad(!src_data_200),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(int_output_sel_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_output_sel[1]~2 .extended_lut = "off";
defparam \int_output_sel[1]~2 .lut_mask = 64'h5303530353035303;
defparam \int_output_sel[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!src_data_198),
	.datab(!src_data_199),
	.datac(!src_data_200),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'h1010101010101010;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \in_ready~1 (
	.dataa(!saved_grant_1),
	.datab(!src_data_198),
	.datac(!src_data_199),
	.datad(!src_data_200),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_ready~1 .extended_lut = "off";
defparam \in_ready~1 .lut_mask = 64'h02AA02AA02AA02AA;
defparam \in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \count~0 (
	.dataa(!\in_ready~1_combout ),
	.datab(!nxt_in_ready),
	.datac(!nxt_in_ready1),
	.datad(!WideOr1),
	.datae(!use_reg1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~0 .extended_lut = "off";
defparam \count~0 .lut_mask = 64'h0051F3F30051F3F3;
defparam \count~0 .shared_arith = "off";

dffeas \count[0] (
	.clk(outclk_wire_0),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count~0_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!src_data_198),
	.datab(!src_data_199),
	.datac(!src_data_200),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'h2020202020202020;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\count[0]~q ),
	.datab(!use_reg1),
	.datac(!\Decoder0~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'hE2E2E2E2E2E2E2E2;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\count[1]~q ),
	.datab(!\Decoder0~0_combout ),
	.datac(!use_reg1),
	.datad(!\Add0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h35CA35CA35CA35CA;
defparam \Add0~1 .shared_arith = "off";

dffeas \count[1] (
	.clk(outclk_wire_0),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count~0_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cyclonev_lcell_comb \out_endofpacket~0 (
	.dataa(!\count[1]~q ),
	.datab(!\count[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_endofpacket~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_endofpacket~0 .extended_lut = "off";
defparam \out_endofpacket~0 .lut_mask = 64'h2222222222222222;
defparam \out_endofpacket~0 .shared_arith = "off";

cyclonev_lcell_comb \use_reg~0 (
	.dataa(!\out_endofpacket~0_combout ),
	.datab(!\in_ready~1_combout ),
	.datac(!nxt_in_ready),
	.datad(!nxt_in_ready1),
	.datae(!WideOr1),
	.dataf(!use_reg1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\use_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \use_reg~0 .extended_lut = "off";
defparam \use_reg~0 .lut_mask = 64'h00003303AAFAAAFA;
defparam \use_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~3 (
	.dataa(!src_data_198),
	.datab(!src_data_199),
	.datac(!src_data_200),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~3 .extended_lut = "off";
defparam \Decoder0~3 .lut_mask = 64'h0202020202020202;
defparam \Decoder0~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~4 (
	.dataa(!src_data_198),
	.datab(!src_data_199),
	.datac(!src_data_200),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~4 .extended_lut = "off";
defparam \Decoder0~4 .lut_mask = 64'h0101010101010101;
defparam \Decoder0~4 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~2 (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_ARSIZE_2),
	.datac(!h2f_AWSIZE_1),
	.datad(!h2f_AWSIZE_2),
	.datae(!saved_grant_1),
	.dataf(!saved_grant_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~2 .extended_lut = "off";
defparam \Decoder0~2 .lut_mask = 64'hFFFF8888F0008000;
defparam \Decoder0~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~5 (
	.dataa(!src_data_198),
	.datab(!\Decoder0~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~5 .extended_lut = "off";
defparam \Decoder0~5 .lut_mask = 64'h1111111111111111;
defparam \Decoder0~5 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~0 (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_ARSIZE_2),
	.datac(!h2f_AWSIZE_1),
	.datad(!h2f_AWSIZE_2),
	.datae(!saved_grant_1),
	.dataf(!saved_grant_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~0 .extended_lut = "off";
defparam \LessThan3~0 .lut_mask = 64'h000066660FF06CA0;
defparam \LessThan3~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~6 (
	.dataa(!src_data_198),
	.datab(!\Decoder0~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~6 .extended_lut = "off";
defparam \Decoder0~6 .lut_mask = 64'h2222222222222222;
defparam \Decoder0~6 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(!\Decoder0~3_combout ),
	.datab(!\Decoder0~4_combout ),
	.datac(!\Decoder0~6_combout ),
	.datad(!out_data_36),
	.datae(gnd),
	.dataf(!\LessThan3~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000F7FF000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\Decoder0~3_combout ),
	.datab(!\Decoder0~4_combout ),
	.datac(!\Decoder0~5_combout ),
	.datad(!out_data_37),
	.datae(gnd),
	.dataf(!\LessThan3~0_combout ),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000F7FF000000FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \address_reg~0 (
	.dataa(!nxt_in_ready),
	.datab(!nxt_in_ready1),
	.datac(!use_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\address_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \address_reg~0 .extended_lut = "off";
defparam \address_reg~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \address_reg~0 .shared_arith = "off";

dffeas \address_reg[1] (
	.clk(outclk_wire_0),
	.d(\Add1~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\address_reg[1]~q ),
	.prn(vcc));
defparam \address_reg[1] .is_wysiwyg = "true";
defparam \address_reg[1] .power_up = "low";

cyclonev_lcell_comb \out_data[37]~2 (
	.dataa(!h2f_ARADDR_1),
	.datab(!h2f_AWADDR_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(!sop_enable),
	.dataf(!address_burst_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[37]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[37]~2 .extended_lut = "off";
defparam \out_data[37]~2 .lut_mask = 64'h05370505053705FF;
defparam \out_data[37]~2 .shared_arith = "off";

dffeas \address_reg[0] (
	.clk(outclk_wire_0),
	.d(\Add1~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\address_reg[0]~q ),
	.prn(vcc));
defparam \address_reg[0] .is_wysiwyg = "true";
defparam \address_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add1~9 (
	.dataa(!\LessThan3~0_combout ),
	.datab(!\Decoder0~3_combout ),
	.datac(!\Decoder0~4_combout ),
	.datad(!int_output_sel_0),
	.datae(gnd),
	.dataf(!\Decoder0~1_combout ),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h00008000000000FF;
defparam \Add1~9 .shared_arith = "off";

dffeas \address_reg[2] (
	.clk(outclk_wire_0),
	.d(\Add1~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\address_reg[2]~q ),
	.prn(vcc));
defparam \address_reg[2] .is_wysiwyg = "true";
defparam \address_reg[2] .power_up = "low";

dffeas endofpacket_reg(
	.clk(outclk_wire_0),
	.d(in_endofpacket),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!use_reg1),
	.q(\endofpacket_reg~q ),
	.prn(vcc));
defparam endofpacket_reg.is_wysiwyg = "true";
defparam endofpacket_reg.power_up = "low";

cyclonev_lcell_comb \LessThan2~0 (
	.dataa(!src_data_198),
	.datab(!src_data_199),
	.datac(!src_data_200),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~0 .extended_lut = "off";
defparam \LessThan2~0 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \LessThan2~0 .shared_arith = "off";

cyclonev_lcell_comb \out_endofpacket~1 (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(!\LessThan2~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_endofpacket~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_endofpacket~1 .extended_lut = "off";
defparam \out_endofpacket~1 .lut_mask = 64'hCCC8CCC8CCC8CCC8;
defparam \out_endofpacket~1 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~6 (
	.dataa(!src_data_198),
	.datab(!src_data_199),
	.datac(!src_data_200),
	.datad(!src_data_184),
	.datae(!src_data_186),
	.dataf(!src_data_185),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~6 .extended_lut = "off";
defparam \ShiftLeft0~6 .lut_mask = 64'h00E208EA04E60CEE;
defparam \ShiftLeft0~6 .shared_arith = "off";

cyclonev_lcell_comb \byte_cnt_reg~0 (
	.dataa(!src_data_200),
	.datab(!nxt_in_ready),
	.datac(!nxt_in_ready1),
	.datad(!use_reg1),
	.datae(!\byte_cnt_reg[2]~q ),
	.dataf(!\ShiftLeft0~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\byte_cnt_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \byte_cnt_reg~0 .extended_lut = "off";
defparam \byte_cnt_reg~0 .lut_mask = 64'hFFF3FF0C55F3550C;
defparam \byte_cnt_reg~0 .shared_arith = "off";

dffeas \byte_cnt_reg[2] (
	.clk(outclk_wire_0),
	.d(\byte_cnt_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byte_cnt_reg[2]~q ),
	.prn(vcc));
defparam \byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \byte_cnt_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!src_data_198),
	.datab(!\Decoder0~2_combout ),
	.datac(!src_data_184),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h0B0B0B0B0B0B0B0B;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \int_byte_cnt_factor[0]~0 (
	.dataa(!src_data_198),
	.datab(!\Decoder0~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_byte_cnt_factor[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_byte_cnt_factor[0]~0 .extended_lut = "off";
defparam \int_byte_cnt_factor[0]~0 .lut_mask = 64'h4444444444444444;
defparam \int_byte_cnt_factor[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_ARSIZE_2),
	.datac(!h2f_AWSIZE_1),
	.datad(!h2f_AWSIZE_2),
	.datae(!saved_grant_1),
	.dataf(!saved_grant_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h0000222200F020A0;
defparam \ShiftLeft0~2 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!src_data_187),
	.datab(!src_data_186),
	.datac(!src_data_185),
	.datad(!src_data_184),
	.datae(!\int_byte_cnt_factor[0]~0_combout ),
	.dataf(!\ShiftLeft0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'h0F0F00FF55553333;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~7 (
	.dataa(!src_data_200),
	.datab(!\Decoder0~0_combout ),
	.datac(!\ShiftLeft0~3_combout ),
	.datad(!src_data_188),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~7 .extended_lut = "off";
defparam \ShiftLeft0~7 .lut_mask = 64'h3705370537053705;
defparam \ShiftLeft0~7 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!src_data_198),
	.datab(!\Decoder0~2_combout ),
	.datac(!src_payload),
	.datad(!src_payload1),
	.datae(!src_payload2),
	.dataf(!src_payload3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'hF444B000B000B000;
defparam \ShiftLeft0~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[78]~12 (
	.dataa(!saved_grant_0),
	.datab(!src_data_198),
	.datac(!\Decoder0~2_combout ),
	.datad(!write_cp_data_187),
	.datae(!src_payload5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[78]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[78]~12 .extended_lut = "off";
defparam \out_data[78]~12 .lut_mask = 64'h0010303000103030;
defparam \out_data[78]~12 .shared_arith = "off";

cyclonev_lcell_comb \out_data[78]~13 (
	.dataa(!saved_grant_0),
	.datab(!src_data_198),
	.datac(!\Decoder0~2_combout ),
	.datad(!write_cp_data_188),
	.datae(!src_payload4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[78]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[78]~13 .extended_lut = "off";
defparam \out_data[78]~13 .lut_mask = 64'h0045CFCF0045CFCF;
defparam \out_data[78]~13 .shared_arith = "off";

cyclonev_lcell_comb \out_data[78]~20 (
	.dataa(!src_data_199),
	.datab(!src_data_200),
	.datac(!\ShiftLeft0~0_combout ),
	.datad(!\ShiftLeft0~1_combout ),
	.datae(!\out_data[78]~12_combout ),
	.dataf(!\out_data[78]~13_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[78]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[78]~20 .extended_lut = "off";
defparam \out_data[78]~20 .lut_mask = 64'h2301EFCDEFCDEFCD;
defparam \out_data[78]~20 .shared_arith = "off";

cyclonev_lcell_comb \out_data[77]~8 (
	.dataa(!src_data_198),
	.datab(!src_data_199),
	.datac(!src_data_200),
	.datad(!src_data_184),
	.datae(!src_payload2),
	.dataf(!src_payload3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[77]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[77]~8 .extended_lut = "off";
defparam \out_data[77]~8 .lut_mask = 64'h0004080C080C080C;
defparam \out_data[77]~8 .shared_arith = "off";

cyclonev_lcell_comb \out_data[77]~9 (
	.dataa(!src_data_198),
	.datab(!\Decoder0~2_combout ),
	.datac(!src_payload),
	.datad(!src_payload1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[77]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[77]~9 .extended_lut = "off";
defparam \out_data[77]~9 .lut_mask = 64'h0444044404440444;
defparam \out_data[77]~9 .shared_arith = "off";

cyclonev_lcell_comb \out_data[77]~10 (
	.dataa(!saved_grant_0),
	.datab(!src_data_198),
	.datac(!\Decoder0~2_combout ),
	.datad(!write_cp_data_187),
	.datae(!src_payload5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[77]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[77]~10 .extended_lut = "off";
defparam \out_data[77]~10 .lut_mask = 64'h0045CFCF0045CFCF;
defparam \out_data[77]~10 .shared_arith = "off";

cyclonev_lcell_comb \out_data[77]~19 (
	.dataa(!src_data_200),
	.datab(!\out_data[77]~8_combout ),
	.datac(!\out_data[77]~9_combout ),
	.datad(!\out_data[77]~10_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[77]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[77]~19 .extended_lut = "off";
defparam \out_data[77]~19 .lut_mask = 64'h3BBB3BBB3BBB3BBB;
defparam \out_data[77]~19 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!src_data_198),
	.datab(!src_data_199),
	.datac(!src_data_200),
	.datad(!src_data_184),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h0008000800080008;
defparam \ShiftLeft0~4 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~5 (
	.dataa(!src_data_188),
	.datab(!src_data_187),
	.datac(!src_data_186),
	.datad(!src_data_185),
	.datae(!\int_byte_cnt_factor[0]~0_combout ),
	.dataf(!\ShiftLeft0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~5 .extended_lut = "off";
defparam \ShiftLeft0~5 .lut_mask = 64'h0F0F00FFAAAA3333;
defparam \ShiftLeft0~5 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~8 (
	.dataa(!src_data_200),
	.datab(!\ShiftLeft0~4_combout ),
	.datac(!\ShiftLeft0~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~8 .extended_lut = "off";
defparam \ShiftLeft0~8 .lut_mask = 64'h3B3B3B3B3B3B3B3B;
defparam \ShiftLeft0~8 .shared_arith = "off";

cyclonev_lcell_comb \Add2~26 (
	.dataa(!use_reg1),
	.datab(!src_data_200),
	.datac(!\byte_cnt_reg[2]~q ),
	.datad(!\ShiftLeft0~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add2~26_cout ),
	.shareout());
defparam \Add2~26 .extended_lut = "off";
defparam \Add2~26 .lut_mask = 64'h000000000000058D;
defparam \Add2~26 .shared_arith = "off";

cyclonev_lcell_comb \Add2~21 (
	.dataa(!use_reg1),
	.datab(!src_data_200),
	.datac(!\ShiftLeft0~3_combout ),
	.datad(!\byte_cnt_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~26_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~21_sumout ),
	.cout(\Add2~22 ),
	.shareout());
defparam \Add2~21 .extended_lut = "off";
defparam \Add2~21 .lut_mask = 64'h000000000000085D;
defparam \Add2~21 .shared_arith = "off";

dffeas \byte_cnt_reg[3] (
	.clk(outclk_wire_0),
	.d(\Add2~21_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\byte_cnt_reg[3]~q ),
	.prn(vcc));
defparam \byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \byte_cnt_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add2~5 (
	.dataa(!use_reg1),
	.datab(gnd),
	.datac(!\byte_cnt_reg[4]~q ),
	.datad(!\ShiftLeft0~8_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h00000000000005AF;
defparam \Add2~5 .shared_arith = "off";

dffeas \byte_cnt_reg[4] (
	.clk(outclk_wire_0),
	.d(\Add2~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\byte_cnt_reg[4]~q ),
	.prn(vcc));
defparam \byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \byte_cnt_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add2~9 (
	.dataa(!use_reg1),
	.datab(gnd),
	.datac(!\byte_cnt_reg[5]~q ),
	.datad(!\out_data[77]~19_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h00000000000005AF;
defparam \Add2~9 .shared_arith = "off";

dffeas \byte_cnt_reg[5] (
	.clk(outclk_wire_0),
	.d(\Add2~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\byte_cnt_reg[5]~q ),
	.prn(vcc));
defparam \byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \byte_cnt_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add2~13 (
	.dataa(!use_reg1),
	.datab(gnd),
	.datac(!\byte_cnt_reg[6]~q ),
	.datad(!\out_data[78]~20_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h00000000000005AF;
defparam \Add2~13 .shared_arith = "off";

dffeas \byte_cnt_reg[6] (
	.clk(outclk_wire_0),
	.d(\Add2~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\byte_cnt_reg[6]~q ),
	.prn(vcc));
defparam \byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \byte_cnt_reg[6] .power_up = "low";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!use_reg1),
	.datab(gnd),
	.datac(!\byte_cnt_reg[7]~q ),
	.datad(!\ShiftLeft0~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h00000000000005AF;
defparam \Add2~1 .shared_arith = "off";

dffeas \byte_cnt_reg[7] (
	.clk(outclk_wire_0),
	.d(\Add2~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\byte_cnt_reg[7]~q ),
	.prn(vcc));
defparam \byte_cnt_reg[7] .is_wysiwyg = "true";
defparam \byte_cnt_reg[7] .power_up = "low";

cyclonev_lcell_comb \Add2~17 (
	.dataa(!use_reg1),
	.datab(!src_data_200),
	.datac(!\ShiftLeft0~5_combout ),
	.datad(!\byte_cnt_reg[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~17_sumout ),
	.cout(),
	.shareout());
defparam \Add2~17 .extended_lut = "off";
defparam \Add2~17 .lut_mask = 64'h0000000000000257;
defparam \Add2~17 .shared_arith = "off";

dffeas \byte_cnt_reg[8] (
	.clk(outclk_wire_0),
	.d(\Add2~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\byte_cnt_reg[8]~q ),
	.prn(vcc));
defparam \byte_cnt_reg[8] .is_wysiwyg = "true";
defparam \byte_cnt_reg[8] .power_up = "low";

cyclonev_lcell_comb \Add1~13 (
	.dataa(!\LessThan3~0_combout ),
	.datab(!\Decoder0~3_combout ),
	.datac(!\Decoder0~4_combout ),
	.datad(!int_output_sel_1),
	.datae(gnd),
	.dataf(!\Decoder0~0_combout ),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FF7F000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(!saved_grant_0),
	.datab(!use_reg1),
	.datac(!out_data_4),
	.datad(!src_payload6),
	.datae(gnd),
	.dataf(!address_reg_4),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFCC000004CC;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(!saved_grant_0),
	.datab(!use_reg1),
	.datac(!out_data_5),
	.datad(!src_payload7),
	.datae(gnd),
	.dataf(!address_reg_5),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFCC000004CC;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(!saved_grant_0),
	.datab(!use_reg1),
	.datac(!out_data_6),
	.datad(!src_payload8),
	.datae(gnd),
	.dataf(!address_reg_6),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h0000FFCC000004CC;
defparam \Add1~25 .shared_arith = "off";

cyclonev_lcell_comb \Add1~29 (
	.dataa(!saved_grant_0),
	.datab(!use_reg1),
	.datac(!out_data_7),
	.datad(!src_payload9),
	.datae(gnd),
	.dataf(!address_reg_7),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~29_sumout ),
	.cout(\Add1~30 ),
	.shareout());
defparam \Add1~29 .extended_lut = "off";
defparam \Add1~29 .lut_mask = 64'h0000FFCC000004CC;
defparam \Add1~29 .shared_arith = "off";

cyclonev_lcell_comb \Add1~33 (
	.dataa(!use_reg1),
	.datab(gnd),
	.datac(!\address_reg[8]~q ),
	.datad(!src_data_152),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~33_sumout ),
	.cout(\Add1~34 ),
	.shareout());
defparam \Add1~33 .extended_lut = "off";
defparam \Add1~33 .lut_mask = 64'h0000FFFF000005AF;
defparam \Add1~33 .shared_arith = "off";

dffeas \address_reg[8] (
	.clk(outclk_wire_0),
	.d(\Add1~33_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\address_reg[8]~q ),
	.prn(vcc));
defparam \address_reg[8] .is_wysiwyg = "true";
defparam \address_reg[8] .power_up = "low";

cyclonev_lcell_comb \Add1~37 (
	.dataa(!use_reg1),
	.datab(!src_payload11),
	.datac(!\address_reg[9]~q ),
	.datad(!src_payload10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~37_sumout ),
	.cout(),
	.shareout());
defparam \Add1~37 .extended_lut = "off";
defparam \Add1~37 .lut_mask = 64'h0000FFFF000027AF;
defparam \Add1~37 .shared_arith = "off";

dffeas \address_reg[9] (
	.clk(outclk_wire_0),
	.d(\Add1~37_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\address_reg[9]~q ),
	.prn(vcc));
defparam \address_reg[9] .is_wysiwyg = "true";
defparam \address_reg[9] .power_up = "low";

cyclonev_lcell_comb \int_output_sel[1]~1 (
	.dataa(!h2f_ARADDR_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(!out_data_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_output_sel[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_output_sel[1]~1 .extended_lut = "off";
defparam \int_output_sel[1]~1 .lut_mask = 64'h111F111F111F111F;
defparam \int_output_sel[1]~1 .shared_arith = "off";

dffeas \address_reg[3] (
	.clk(outclk_wire_0),
	.d(\Add1~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address_reg~0_combout ),
	.q(\address_reg[3]~q ),
	.prn(vcc));
defparam \address_reg[3] .is_wysiwyg = "true";
defparam \address_reg[3] .power_up = "low";

endmodule

module Computer_System_altera_merlin_width_adapter_3 (
	h2f_BREADY_0,
	h2f_RREADY_0,
	q_b_0,
	q_b_2,
	q_b_3,
	q_b_5,
	q_b_7,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_18,
	q_b_19,
	q_b_21,
	q_b_23,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_30,
	q_b_31,
	outclk_wire_0,
	data_reg_0,
	data_reg_1,
	data_reg_2,
	data_reg_3,
	data_reg_4,
	data_reg_5,
	data_reg_6,
	data_reg_7,
	data_reg_8,
	data_reg_9,
	data_reg_10,
	data_reg_11,
	data_reg_12,
	data_reg_13,
	data_reg_14,
	data_reg_15,
	data_reg_16,
	data_reg_17,
	data_reg_18,
	data_reg_19,
	data_reg_20,
	data_reg_21,
	data_reg_22,
	data_reg_23,
	data_reg_24,
	data_reg_25,
	data_reg_26,
	data_reg_27,
	data_reg_28,
	data_reg_29,
	data_reg_30,
	data_reg_31,
	data_reg_32,
	data_reg_33,
	data_reg_34,
	data_reg_35,
	data_reg_36,
	data_reg_37,
	data_reg_38,
	data_reg_39,
	data_reg_40,
	data_reg_41,
	data_reg_42,
	data_reg_43,
	data_reg_44,
	data_reg_45,
	data_reg_46,
	data_reg_47,
	data_reg_48,
	data_reg_49,
	data_reg_50,
	data_reg_51,
	data_reg_52,
	data_reg_53,
	data_reg_54,
	data_reg_55,
	data_reg_56,
	data_reg_57,
	data_reg_58,
	data_reg_59,
	data_reg_60,
	data_reg_61,
	data_reg_62,
	data_reg_63,
	data_reg_64,
	data_reg_65,
	data_reg_66,
	data_reg_67,
	data_reg_68,
	data_reg_69,
	data_reg_70,
	data_reg_71,
	data_reg_72,
	data_reg_73,
	data_reg_74,
	data_reg_75,
	data_reg_76,
	data_reg_77,
	data_reg_78,
	data_reg_79,
	data_reg_80,
	data_reg_81,
	data_reg_82,
	data_reg_83,
	data_reg_84,
	data_reg_85,
	data_reg_86,
	data_reg_87,
	data_reg_88,
	data_reg_89,
	data_reg_90,
	data_reg_91,
	data_reg_92,
	data_reg_93,
	data_reg_94,
	data_reg_95,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_125_0,
	mem_used_01,
	out_valid,
	comb,
	burst_uncompress_busy,
	src_payload,
	mem_38_0,
	source_addr_2,
	source_addr_21,
	mem_122_0,
	mem_123_0,
	mem_91_0,
	mem_124_0,
	mem_90_0,
	mem_39_0,
	source_addr_3,
	always10,
	src0_valid,
	ShiftLeft0,
	always4,
	mem_0_0,
	LessThan15,
	mem_2_0,
	mem_3_0,
	mem_5_0,
	mem_7_0,
	mem_9_0,
	mem_10_0,
	mem_11_0,
	mem_12_0,
	mem_14_0,
	mem_15_0,
	mem_16_0,
	mem_18_0,
	mem_19_0,
	mem_21_0,
	mem_23_0,
	mem_25_0,
	mem_26_0,
	mem_27_0,
	mem_28_0,
	mem_30_0,
	mem_31_0,
	ShiftLeft01,
	ShiftLeft02,
	out_data_1,
	out_data_4,
	out_data_6,
	out_data_8,
	out_data_13,
	out_data_17,
	out_data_20,
	out_data_22,
	out_data_24,
	out_data_29,
	r_sync_rst,
	p1_ready,
	always101)/* synthesis synthesis_greybox=0 */;
input 	h2f_BREADY_0;
input 	h2f_RREADY_0;
input 	q_b_0;
input 	q_b_2;
input 	q_b_3;
input 	q_b_5;
input 	q_b_7;
input 	q_b_9;
input 	q_b_10;
input 	q_b_11;
input 	q_b_12;
input 	q_b_14;
input 	q_b_15;
input 	q_b_16;
input 	q_b_18;
input 	q_b_19;
input 	q_b_21;
input 	q_b_23;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_28;
input 	q_b_30;
input 	q_b_31;
input 	outclk_wire_0;
output 	data_reg_0;
output 	data_reg_1;
output 	data_reg_2;
output 	data_reg_3;
output 	data_reg_4;
output 	data_reg_5;
output 	data_reg_6;
output 	data_reg_7;
output 	data_reg_8;
output 	data_reg_9;
output 	data_reg_10;
output 	data_reg_11;
output 	data_reg_12;
output 	data_reg_13;
output 	data_reg_14;
output 	data_reg_15;
output 	data_reg_16;
output 	data_reg_17;
output 	data_reg_18;
output 	data_reg_19;
output 	data_reg_20;
output 	data_reg_21;
output 	data_reg_22;
output 	data_reg_23;
output 	data_reg_24;
output 	data_reg_25;
output 	data_reg_26;
output 	data_reg_27;
output 	data_reg_28;
output 	data_reg_29;
output 	data_reg_30;
output 	data_reg_31;
output 	data_reg_32;
output 	data_reg_33;
output 	data_reg_34;
output 	data_reg_35;
output 	data_reg_36;
output 	data_reg_37;
output 	data_reg_38;
output 	data_reg_39;
output 	data_reg_40;
output 	data_reg_41;
output 	data_reg_42;
output 	data_reg_43;
output 	data_reg_44;
output 	data_reg_45;
output 	data_reg_46;
output 	data_reg_47;
output 	data_reg_48;
output 	data_reg_49;
output 	data_reg_50;
output 	data_reg_51;
output 	data_reg_52;
output 	data_reg_53;
output 	data_reg_54;
output 	data_reg_55;
output 	data_reg_56;
output 	data_reg_57;
output 	data_reg_58;
output 	data_reg_59;
output 	data_reg_60;
output 	data_reg_61;
output 	data_reg_62;
output 	data_reg_63;
output 	data_reg_64;
output 	data_reg_65;
output 	data_reg_66;
output 	data_reg_67;
output 	data_reg_68;
output 	data_reg_69;
output 	data_reg_70;
output 	data_reg_71;
output 	data_reg_72;
output 	data_reg_73;
output 	data_reg_74;
output 	data_reg_75;
output 	data_reg_76;
output 	data_reg_77;
output 	data_reg_78;
output 	data_reg_79;
output 	data_reg_80;
output 	data_reg_81;
output 	data_reg_82;
output 	data_reg_83;
output 	data_reg_84;
output 	data_reg_85;
output 	data_reg_86;
output 	data_reg_87;
output 	data_reg_88;
output 	data_reg_89;
output 	data_reg_90;
output 	data_reg_91;
output 	data_reg_92;
output 	data_reg_93;
output 	data_reg_94;
output 	data_reg_95;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_125_0;
input 	mem_used_01;
output 	out_valid;
input 	comb;
input 	burst_uncompress_busy;
input 	src_payload;
input 	mem_38_0;
input 	source_addr_2;
input 	source_addr_21;
input 	mem_122_0;
input 	mem_123_0;
input 	mem_91_0;
input 	mem_124_0;
input 	mem_90_0;
input 	mem_39_0;
input 	source_addr_3;
output 	always10;
input 	src0_valid;
output 	ShiftLeft0;
input 	always4;
input 	mem_0_0;
output 	LessThan15;
input 	mem_2_0;
input 	mem_3_0;
input 	mem_5_0;
input 	mem_7_0;
input 	mem_9_0;
input 	mem_10_0;
input 	mem_11_0;
input 	mem_12_0;
input 	mem_14_0;
input 	mem_15_0;
input 	mem_16_0;
input 	mem_18_0;
input 	mem_19_0;
input 	mem_21_0;
input 	mem_23_0;
input 	mem_25_0;
input 	mem_26_0;
input 	mem_27_0;
input 	mem_28_0;
input 	mem_30_0;
input 	mem_31_0;
output 	ShiftLeft01;
output 	ShiftLeft02;
input 	out_data_1;
input 	out_data_4;
input 	out_data_6;
input 	out_data_8;
input 	out_data_13;
input 	out_data_17;
input 	out_data_20;
input 	out_data_22;
input 	out_data_24;
input 	out_data_29;
input 	r_sync_rst;
output 	p1_ready;
output 	always101;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_reg~0_combout ;
wire \always9~0_combout ;
wire \data_reg~1_combout ;
wire \data_reg~2_combout ;
wire \data_reg~3_combout ;
wire \data_reg~4_combout ;
wire \data_reg~5_combout ;
wire \data_reg~6_combout ;
wire \data_reg~7_combout ;
wire \data_reg~8_combout ;
wire \data_reg~9_combout ;
wire \data_reg~10_combout ;
wire \data_reg~11_combout ;
wire \data_reg~12_combout ;
wire \data_reg~13_combout ;
wire \data_reg~14_combout ;
wire \data_reg~15_combout ;
wire \data_reg~16_combout ;
wire \data_reg~17_combout ;
wire \data_reg~18_combout ;
wire \data_reg~19_combout ;
wire \data_reg~20_combout ;
wire \data_reg~21_combout ;
wire \data_reg~22_combout ;
wire \data_reg~23_combout ;
wire \data_reg~24_combout ;
wire \data_reg~25_combout ;
wire \data_reg~26_combout ;
wire \data_reg~27_combout ;
wire \data_reg~28_combout ;
wire \data_reg~29_combout ;
wire \data_reg~30_combout ;
wire \data_reg~31_combout ;
wire \data_reg~32_combout ;
wire \data_reg~33_combout ;
wire \data_reg~34_combout ;
wire \data_reg~35_combout ;
wire \data_reg~36_combout ;
wire \data_reg~37_combout ;
wire \data_reg~38_combout ;
wire \data_reg~39_combout ;
wire \data_reg~40_combout ;
wire \data_reg~41_combout ;
wire \data_reg~42_combout ;
wire \data_reg~43_combout ;
wire \data_reg~44_combout ;
wire \data_reg~45_combout ;
wire \data_reg~46_combout ;
wire \data_reg~47_combout ;
wire \data_reg~48_combout ;
wire \data_reg~49_combout ;
wire \data_reg~50_combout ;
wire \data_reg~51_combout ;
wire \data_reg~52_combout ;
wire \data_reg~53_combout ;
wire \data_reg~54_combout ;
wire \data_reg~55_combout ;
wire \data_reg~56_combout ;
wire \data_reg~57_combout ;
wire \data_reg~58_combout ;
wire \data_reg~59_combout ;
wire \data_reg~60_combout ;
wire \data_reg~61_combout ;
wire \data_reg~62_combout ;
wire \data_reg~63_combout ;
wire \data_reg~64_combout ;
wire \data_reg~65_combout ;
wire \data_reg~66_combout ;
wire \data_reg~67_combout ;
wire \data_reg~68_combout ;
wire \data_reg~69_combout ;
wire \data_reg~70_combout ;
wire \data_reg~71_combout ;
wire \data_reg~72_combout ;
wire \data_reg~73_combout ;
wire \data_reg~74_combout ;
wire \data_reg~75_combout ;
wire \data_reg~76_combout ;
wire \data_reg~77_combout ;
wire \data_reg~78_combout ;
wire \data_reg~79_combout ;
wire \data_reg~80_combout ;
wire \data_reg~81_combout ;
wire \data_reg~82_combout ;
wire \data_reg~83_combout ;
wire \data_reg~84_combout ;
wire \data_reg~85_combout ;
wire \data_reg~86_combout ;
wire \data_reg~87_combout ;
wire \data_reg~88_combout ;
wire \data_reg~89_combout ;
wire \data_reg~90_combout ;
wire \data_reg~91_combout ;
wire \data_reg~92_combout ;
wire \data_reg~93_combout ;
wire \data_reg~94_combout ;
wire \data_reg~95_combout ;
wire \always10~0_combout ;
wire \always10~1_combout ;
wire \ShiftRight0~0_combout ;
wire \always10~2_combout ;
wire \always10~3_combout ;
wire \always10~4_combout ;
wire \always10~5_combout ;
wire \always10~6_combout ;
wire \always10~7_combout ;
wire \always10~8_combout ;


dffeas \data_reg[0] (
	.clk(outclk_wire_0),
	.d(\data_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_0),
	.prn(vcc));
defparam \data_reg[0] .is_wysiwyg = "true";
defparam \data_reg[0] .power_up = "low";

dffeas \data_reg[1] (
	.clk(outclk_wire_0),
	.d(\data_reg~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_1),
	.prn(vcc));
defparam \data_reg[1] .is_wysiwyg = "true";
defparam \data_reg[1] .power_up = "low";

dffeas \data_reg[2] (
	.clk(outclk_wire_0),
	.d(\data_reg~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_2),
	.prn(vcc));
defparam \data_reg[2] .is_wysiwyg = "true";
defparam \data_reg[2] .power_up = "low";

dffeas \data_reg[3] (
	.clk(outclk_wire_0),
	.d(\data_reg~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_3),
	.prn(vcc));
defparam \data_reg[3] .is_wysiwyg = "true";
defparam \data_reg[3] .power_up = "low";

dffeas \data_reg[4] (
	.clk(outclk_wire_0),
	.d(\data_reg~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_4),
	.prn(vcc));
defparam \data_reg[4] .is_wysiwyg = "true";
defparam \data_reg[4] .power_up = "low";

dffeas \data_reg[5] (
	.clk(outclk_wire_0),
	.d(\data_reg~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_5),
	.prn(vcc));
defparam \data_reg[5] .is_wysiwyg = "true";
defparam \data_reg[5] .power_up = "low";

dffeas \data_reg[6] (
	.clk(outclk_wire_0),
	.d(\data_reg~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_6),
	.prn(vcc));
defparam \data_reg[6] .is_wysiwyg = "true";
defparam \data_reg[6] .power_up = "low";

dffeas \data_reg[7] (
	.clk(outclk_wire_0),
	.d(\data_reg~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_7),
	.prn(vcc));
defparam \data_reg[7] .is_wysiwyg = "true";
defparam \data_reg[7] .power_up = "low";

dffeas \data_reg[8] (
	.clk(outclk_wire_0),
	.d(\data_reg~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_8),
	.prn(vcc));
defparam \data_reg[8] .is_wysiwyg = "true";
defparam \data_reg[8] .power_up = "low";

dffeas \data_reg[9] (
	.clk(outclk_wire_0),
	.d(\data_reg~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_9),
	.prn(vcc));
defparam \data_reg[9] .is_wysiwyg = "true";
defparam \data_reg[9] .power_up = "low";

dffeas \data_reg[10] (
	.clk(outclk_wire_0),
	.d(\data_reg~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_10),
	.prn(vcc));
defparam \data_reg[10] .is_wysiwyg = "true";
defparam \data_reg[10] .power_up = "low";

dffeas \data_reg[11] (
	.clk(outclk_wire_0),
	.d(\data_reg~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_11),
	.prn(vcc));
defparam \data_reg[11] .is_wysiwyg = "true";
defparam \data_reg[11] .power_up = "low";

dffeas \data_reg[12] (
	.clk(outclk_wire_0),
	.d(\data_reg~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_12),
	.prn(vcc));
defparam \data_reg[12] .is_wysiwyg = "true";
defparam \data_reg[12] .power_up = "low";

dffeas \data_reg[13] (
	.clk(outclk_wire_0),
	.d(\data_reg~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_13),
	.prn(vcc));
defparam \data_reg[13] .is_wysiwyg = "true";
defparam \data_reg[13] .power_up = "low";

dffeas \data_reg[14] (
	.clk(outclk_wire_0),
	.d(\data_reg~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_14),
	.prn(vcc));
defparam \data_reg[14] .is_wysiwyg = "true";
defparam \data_reg[14] .power_up = "low";

dffeas \data_reg[15] (
	.clk(outclk_wire_0),
	.d(\data_reg~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_15),
	.prn(vcc));
defparam \data_reg[15] .is_wysiwyg = "true";
defparam \data_reg[15] .power_up = "low";

dffeas \data_reg[16] (
	.clk(outclk_wire_0),
	.d(\data_reg~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_16),
	.prn(vcc));
defparam \data_reg[16] .is_wysiwyg = "true";
defparam \data_reg[16] .power_up = "low";

dffeas \data_reg[17] (
	.clk(outclk_wire_0),
	.d(\data_reg~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_17),
	.prn(vcc));
defparam \data_reg[17] .is_wysiwyg = "true";
defparam \data_reg[17] .power_up = "low";

dffeas \data_reg[18] (
	.clk(outclk_wire_0),
	.d(\data_reg~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_18),
	.prn(vcc));
defparam \data_reg[18] .is_wysiwyg = "true";
defparam \data_reg[18] .power_up = "low";

dffeas \data_reg[19] (
	.clk(outclk_wire_0),
	.d(\data_reg~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_19),
	.prn(vcc));
defparam \data_reg[19] .is_wysiwyg = "true";
defparam \data_reg[19] .power_up = "low";

dffeas \data_reg[20] (
	.clk(outclk_wire_0),
	.d(\data_reg~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_20),
	.prn(vcc));
defparam \data_reg[20] .is_wysiwyg = "true";
defparam \data_reg[20] .power_up = "low";

dffeas \data_reg[21] (
	.clk(outclk_wire_0),
	.d(\data_reg~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_21),
	.prn(vcc));
defparam \data_reg[21] .is_wysiwyg = "true";
defparam \data_reg[21] .power_up = "low";

dffeas \data_reg[22] (
	.clk(outclk_wire_0),
	.d(\data_reg~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_22),
	.prn(vcc));
defparam \data_reg[22] .is_wysiwyg = "true";
defparam \data_reg[22] .power_up = "low";

dffeas \data_reg[23] (
	.clk(outclk_wire_0),
	.d(\data_reg~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_23),
	.prn(vcc));
defparam \data_reg[23] .is_wysiwyg = "true";
defparam \data_reg[23] .power_up = "low";

dffeas \data_reg[24] (
	.clk(outclk_wire_0),
	.d(\data_reg~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_24),
	.prn(vcc));
defparam \data_reg[24] .is_wysiwyg = "true";
defparam \data_reg[24] .power_up = "low";

dffeas \data_reg[25] (
	.clk(outclk_wire_0),
	.d(\data_reg~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_25),
	.prn(vcc));
defparam \data_reg[25] .is_wysiwyg = "true";
defparam \data_reg[25] .power_up = "low";

dffeas \data_reg[26] (
	.clk(outclk_wire_0),
	.d(\data_reg~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_26),
	.prn(vcc));
defparam \data_reg[26] .is_wysiwyg = "true";
defparam \data_reg[26] .power_up = "low";

dffeas \data_reg[27] (
	.clk(outclk_wire_0),
	.d(\data_reg~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_27),
	.prn(vcc));
defparam \data_reg[27] .is_wysiwyg = "true";
defparam \data_reg[27] .power_up = "low";

dffeas \data_reg[28] (
	.clk(outclk_wire_0),
	.d(\data_reg~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_28),
	.prn(vcc));
defparam \data_reg[28] .is_wysiwyg = "true";
defparam \data_reg[28] .power_up = "low";

dffeas \data_reg[29] (
	.clk(outclk_wire_0),
	.d(\data_reg~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_29),
	.prn(vcc));
defparam \data_reg[29] .is_wysiwyg = "true";
defparam \data_reg[29] .power_up = "low";

dffeas \data_reg[30] (
	.clk(outclk_wire_0),
	.d(\data_reg~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_30),
	.prn(vcc));
defparam \data_reg[30] .is_wysiwyg = "true";
defparam \data_reg[30] .power_up = "low";

dffeas \data_reg[31] (
	.clk(outclk_wire_0),
	.d(\data_reg~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_31),
	.prn(vcc));
defparam \data_reg[31] .is_wysiwyg = "true";
defparam \data_reg[31] .power_up = "low";

dffeas \data_reg[32] (
	.clk(outclk_wire_0),
	.d(\data_reg~32_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_32),
	.prn(vcc));
defparam \data_reg[32] .is_wysiwyg = "true";
defparam \data_reg[32] .power_up = "low";

dffeas \data_reg[33] (
	.clk(outclk_wire_0),
	.d(\data_reg~33_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_33),
	.prn(vcc));
defparam \data_reg[33] .is_wysiwyg = "true";
defparam \data_reg[33] .power_up = "low";

dffeas \data_reg[34] (
	.clk(outclk_wire_0),
	.d(\data_reg~34_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_34),
	.prn(vcc));
defparam \data_reg[34] .is_wysiwyg = "true";
defparam \data_reg[34] .power_up = "low";

dffeas \data_reg[35] (
	.clk(outclk_wire_0),
	.d(\data_reg~35_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_35),
	.prn(vcc));
defparam \data_reg[35] .is_wysiwyg = "true";
defparam \data_reg[35] .power_up = "low";

dffeas \data_reg[36] (
	.clk(outclk_wire_0),
	.d(\data_reg~36_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_36),
	.prn(vcc));
defparam \data_reg[36] .is_wysiwyg = "true";
defparam \data_reg[36] .power_up = "low";

dffeas \data_reg[37] (
	.clk(outclk_wire_0),
	.d(\data_reg~37_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_37),
	.prn(vcc));
defparam \data_reg[37] .is_wysiwyg = "true";
defparam \data_reg[37] .power_up = "low";

dffeas \data_reg[38] (
	.clk(outclk_wire_0),
	.d(\data_reg~38_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_38),
	.prn(vcc));
defparam \data_reg[38] .is_wysiwyg = "true";
defparam \data_reg[38] .power_up = "low";

dffeas \data_reg[39] (
	.clk(outclk_wire_0),
	.d(\data_reg~39_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_39),
	.prn(vcc));
defparam \data_reg[39] .is_wysiwyg = "true";
defparam \data_reg[39] .power_up = "low";

dffeas \data_reg[40] (
	.clk(outclk_wire_0),
	.d(\data_reg~40_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_40),
	.prn(vcc));
defparam \data_reg[40] .is_wysiwyg = "true";
defparam \data_reg[40] .power_up = "low";

dffeas \data_reg[41] (
	.clk(outclk_wire_0),
	.d(\data_reg~41_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_41),
	.prn(vcc));
defparam \data_reg[41] .is_wysiwyg = "true";
defparam \data_reg[41] .power_up = "low";

dffeas \data_reg[42] (
	.clk(outclk_wire_0),
	.d(\data_reg~42_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_42),
	.prn(vcc));
defparam \data_reg[42] .is_wysiwyg = "true";
defparam \data_reg[42] .power_up = "low";

dffeas \data_reg[43] (
	.clk(outclk_wire_0),
	.d(\data_reg~43_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_43),
	.prn(vcc));
defparam \data_reg[43] .is_wysiwyg = "true";
defparam \data_reg[43] .power_up = "low";

dffeas \data_reg[44] (
	.clk(outclk_wire_0),
	.d(\data_reg~44_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_44),
	.prn(vcc));
defparam \data_reg[44] .is_wysiwyg = "true";
defparam \data_reg[44] .power_up = "low";

dffeas \data_reg[45] (
	.clk(outclk_wire_0),
	.d(\data_reg~45_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_45),
	.prn(vcc));
defparam \data_reg[45] .is_wysiwyg = "true";
defparam \data_reg[45] .power_up = "low";

dffeas \data_reg[46] (
	.clk(outclk_wire_0),
	.d(\data_reg~46_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_46),
	.prn(vcc));
defparam \data_reg[46] .is_wysiwyg = "true";
defparam \data_reg[46] .power_up = "low";

dffeas \data_reg[47] (
	.clk(outclk_wire_0),
	.d(\data_reg~47_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_47),
	.prn(vcc));
defparam \data_reg[47] .is_wysiwyg = "true";
defparam \data_reg[47] .power_up = "low";

dffeas \data_reg[48] (
	.clk(outclk_wire_0),
	.d(\data_reg~48_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_48),
	.prn(vcc));
defparam \data_reg[48] .is_wysiwyg = "true";
defparam \data_reg[48] .power_up = "low";

dffeas \data_reg[49] (
	.clk(outclk_wire_0),
	.d(\data_reg~49_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_49),
	.prn(vcc));
defparam \data_reg[49] .is_wysiwyg = "true";
defparam \data_reg[49] .power_up = "low";

dffeas \data_reg[50] (
	.clk(outclk_wire_0),
	.d(\data_reg~50_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_50),
	.prn(vcc));
defparam \data_reg[50] .is_wysiwyg = "true";
defparam \data_reg[50] .power_up = "low";

dffeas \data_reg[51] (
	.clk(outclk_wire_0),
	.d(\data_reg~51_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_51),
	.prn(vcc));
defparam \data_reg[51] .is_wysiwyg = "true";
defparam \data_reg[51] .power_up = "low";

dffeas \data_reg[52] (
	.clk(outclk_wire_0),
	.d(\data_reg~52_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_52),
	.prn(vcc));
defparam \data_reg[52] .is_wysiwyg = "true";
defparam \data_reg[52] .power_up = "low";

dffeas \data_reg[53] (
	.clk(outclk_wire_0),
	.d(\data_reg~53_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_53),
	.prn(vcc));
defparam \data_reg[53] .is_wysiwyg = "true";
defparam \data_reg[53] .power_up = "low";

dffeas \data_reg[54] (
	.clk(outclk_wire_0),
	.d(\data_reg~54_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_54),
	.prn(vcc));
defparam \data_reg[54] .is_wysiwyg = "true";
defparam \data_reg[54] .power_up = "low";

dffeas \data_reg[55] (
	.clk(outclk_wire_0),
	.d(\data_reg~55_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_55),
	.prn(vcc));
defparam \data_reg[55] .is_wysiwyg = "true";
defparam \data_reg[55] .power_up = "low";

dffeas \data_reg[56] (
	.clk(outclk_wire_0),
	.d(\data_reg~56_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_56),
	.prn(vcc));
defparam \data_reg[56] .is_wysiwyg = "true";
defparam \data_reg[56] .power_up = "low";

dffeas \data_reg[57] (
	.clk(outclk_wire_0),
	.d(\data_reg~57_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_57),
	.prn(vcc));
defparam \data_reg[57] .is_wysiwyg = "true";
defparam \data_reg[57] .power_up = "low";

dffeas \data_reg[58] (
	.clk(outclk_wire_0),
	.d(\data_reg~58_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_58),
	.prn(vcc));
defparam \data_reg[58] .is_wysiwyg = "true";
defparam \data_reg[58] .power_up = "low";

dffeas \data_reg[59] (
	.clk(outclk_wire_0),
	.d(\data_reg~59_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_59),
	.prn(vcc));
defparam \data_reg[59] .is_wysiwyg = "true";
defparam \data_reg[59] .power_up = "low";

dffeas \data_reg[60] (
	.clk(outclk_wire_0),
	.d(\data_reg~60_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_60),
	.prn(vcc));
defparam \data_reg[60] .is_wysiwyg = "true";
defparam \data_reg[60] .power_up = "low";

dffeas \data_reg[61] (
	.clk(outclk_wire_0),
	.d(\data_reg~61_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_61),
	.prn(vcc));
defparam \data_reg[61] .is_wysiwyg = "true";
defparam \data_reg[61] .power_up = "low";

dffeas \data_reg[62] (
	.clk(outclk_wire_0),
	.d(\data_reg~62_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_62),
	.prn(vcc));
defparam \data_reg[62] .is_wysiwyg = "true";
defparam \data_reg[62] .power_up = "low";

dffeas \data_reg[63] (
	.clk(outclk_wire_0),
	.d(\data_reg~63_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_63),
	.prn(vcc));
defparam \data_reg[63] .is_wysiwyg = "true";
defparam \data_reg[63] .power_up = "low";

dffeas \data_reg[64] (
	.clk(outclk_wire_0),
	.d(\data_reg~64_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_64),
	.prn(vcc));
defparam \data_reg[64] .is_wysiwyg = "true";
defparam \data_reg[64] .power_up = "low";

dffeas \data_reg[65] (
	.clk(outclk_wire_0),
	.d(\data_reg~65_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_65),
	.prn(vcc));
defparam \data_reg[65] .is_wysiwyg = "true";
defparam \data_reg[65] .power_up = "low";

dffeas \data_reg[66] (
	.clk(outclk_wire_0),
	.d(\data_reg~66_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_66),
	.prn(vcc));
defparam \data_reg[66] .is_wysiwyg = "true";
defparam \data_reg[66] .power_up = "low";

dffeas \data_reg[67] (
	.clk(outclk_wire_0),
	.d(\data_reg~67_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_67),
	.prn(vcc));
defparam \data_reg[67] .is_wysiwyg = "true";
defparam \data_reg[67] .power_up = "low";

dffeas \data_reg[68] (
	.clk(outclk_wire_0),
	.d(\data_reg~68_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_68),
	.prn(vcc));
defparam \data_reg[68] .is_wysiwyg = "true";
defparam \data_reg[68] .power_up = "low";

dffeas \data_reg[69] (
	.clk(outclk_wire_0),
	.d(\data_reg~69_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_69),
	.prn(vcc));
defparam \data_reg[69] .is_wysiwyg = "true";
defparam \data_reg[69] .power_up = "low";

dffeas \data_reg[70] (
	.clk(outclk_wire_0),
	.d(\data_reg~70_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_70),
	.prn(vcc));
defparam \data_reg[70] .is_wysiwyg = "true";
defparam \data_reg[70] .power_up = "low";

dffeas \data_reg[71] (
	.clk(outclk_wire_0),
	.d(\data_reg~71_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_71),
	.prn(vcc));
defparam \data_reg[71] .is_wysiwyg = "true";
defparam \data_reg[71] .power_up = "low";

dffeas \data_reg[72] (
	.clk(outclk_wire_0),
	.d(\data_reg~72_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_72),
	.prn(vcc));
defparam \data_reg[72] .is_wysiwyg = "true";
defparam \data_reg[72] .power_up = "low";

dffeas \data_reg[73] (
	.clk(outclk_wire_0),
	.d(\data_reg~73_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_73),
	.prn(vcc));
defparam \data_reg[73] .is_wysiwyg = "true";
defparam \data_reg[73] .power_up = "low";

dffeas \data_reg[74] (
	.clk(outclk_wire_0),
	.d(\data_reg~74_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_74),
	.prn(vcc));
defparam \data_reg[74] .is_wysiwyg = "true";
defparam \data_reg[74] .power_up = "low";

dffeas \data_reg[75] (
	.clk(outclk_wire_0),
	.d(\data_reg~75_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_75),
	.prn(vcc));
defparam \data_reg[75] .is_wysiwyg = "true";
defparam \data_reg[75] .power_up = "low";

dffeas \data_reg[76] (
	.clk(outclk_wire_0),
	.d(\data_reg~76_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_76),
	.prn(vcc));
defparam \data_reg[76] .is_wysiwyg = "true";
defparam \data_reg[76] .power_up = "low";

dffeas \data_reg[77] (
	.clk(outclk_wire_0),
	.d(\data_reg~77_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_77),
	.prn(vcc));
defparam \data_reg[77] .is_wysiwyg = "true";
defparam \data_reg[77] .power_up = "low";

dffeas \data_reg[78] (
	.clk(outclk_wire_0),
	.d(\data_reg~78_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_78),
	.prn(vcc));
defparam \data_reg[78] .is_wysiwyg = "true";
defparam \data_reg[78] .power_up = "low";

dffeas \data_reg[79] (
	.clk(outclk_wire_0),
	.d(\data_reg~79_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_79),
	.prn(vcc));
defparam \data_reg[79] .is_wysiwyg = "true";
defparam \data_reg[79] .power_up = "low";

dffeas \data_reg[80] (
	.clk(outclk_wire_0),
	.d(\data_reg~80_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_80),
	.prn(vcc));
defparam \data_reg[80] .is_wysiwyg = "true";
defparam \data_reg[80] .power_up = "low";

dffeas \data_reg[81] (
	.clk(outclk_wire_0),
	.d(\data_reg~81_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_81),
	.prn(vcc));
defparam \data_reg[81] .is_wysiwyg = "true";
defparam \data_reg[81] .power_up = "low";

dffeas \data_reg[82] (
	.clk(outclk_wire_0),
	.d(\data_reg~82_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_82),
	.prn(vcc));
defparam \data_reg[82] .is_wysiwyg = "true";
defparam \data_reg[82] .power_up = "low";

dffeas \data_reg[83] (
	.clk(outclk_wire_0),
	.d(\data_reg~83_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_83),
	.prn(vcc));
defparam \data_reg[83] .is_wysiwyg = "true";
defparam \data_reg[83] .power_up = "low";

dffeas \data_reg[84] (
	.clk(outclk_wire_0),
	.d(\data_reg~84_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_84),
	.prn(vcc));
defparam \data_reg[84] .is_wysiwyg = "true";
defparam \data_reg[84] .power_up = "low";

dffeas \data_reg[85] (
	.clk(outclk_wire_0),
	.d(\data_reg~85_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_85),
	.prn(vcc));
defparam \data_reg[85] .is_wysiwyg = "true";
defparam \data_reg[85] .power_up = "low";

dffeas \data_reg[86] (
	.clk(outclk_wire_0),
	.d(\data_reg~86_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_86),
	.prn(vcc));
defparam \data_reg[86] .is_wysiwyg = "true";
defparam \data_reg[86] .power_up = "low";

dffeas \data_reg[87] (
	.clk(outclk_wire_0),
	.d(\data_reg~87_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_87),
	.prn(vcc));
defparam \data_reg[87] .is_wysiwyg = "true";
defparam \data_reg[87] .power_up = "low";

dffeas \data_reg[88] (
	.clk(outclk_wire_0),
	.d(\data_reg~88_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_88),
	.prn(vcc));
defparam \data_reg[88] .is_wysiwyg = "true";
defparam \data_reg[88] .power_up = "low";

dffeas \data_reg[89] (
	.clk(outclk_wire_0),
	.d(\data_reg~89_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_89),
	.prn(vcc));
defparam \data_reg[89] .is_wysiwyg = "true";
defparam \data_reg[89] .power_up = "low";

dffeas \data_reg[90] (
	.clk(outclk_wire_0),
	.d(\data_reg~90_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_90),
	.prn(vcc));
defparam \data_reg[90] .is_wysiwyg = "true";
defparam \data_reg[90] .power_up = "low";

dffeas \data_reg[91] (
	.clk(outclk_wire_0),
	.d(\data_reg~91_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_91),
	.prn(vcc));
defparam \data_reg[91] .is_wysiwyg = "true";
defparam \data_reg[91] .power_up = "low";

dffeas \data_reg[92] (
	.clk(outclk_wire_0),
	.d(\data_reg~92_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_92),
	.prn(vcc));
defparam \data_reg[92] .is_wysiwyg = "true";
defparam \data_reg[92] .power_up = "low";

dffeas \data_reg[93] (
	.clk(outclk_wire_0),
	.d(\data_reg~93_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_93),
	.prn(vcc));
defparam \data_reg[93] .is_wysiwyg = "true";
defparam \data_reg[93] .power_up = "low";

dffeas \data_reg[94] (
	.clk(outclk_wire_0),
	.d(\data_reg~94_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_94),
	.prn(vcc));
defparam \data_reg[94] .is_wysiwyg = "true";
defparam \data_reg[94] .power_up = "low";

dffeas \data_reg[95] (
	.clk(outclk_wire_0),
	.d(\data_reg~95_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(always101),
	.sload(gnd),
	.ena(\always9~0_combout ),
	.q(data_reg_95),
	.prn(vcc));
defparam \data_reg[95] .is_wysiwyg = "true";
defparam \data_reg[95] .power_up = "low";

cyclonev_lcell_comb \out_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_125_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_valid~0 .extended_lut = "off";
defparam \out_valid~0 .lut_mask = 64'h8880888088808880;
defparam \out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \always10~9 (
	.dataa(!source_addr_21),
	.datab(!\always10~1_combout ),
	.datac(!\always10~3_combout ),
	.datad(!\always10~6_combout ),
	.datae(!\always10~7_combout ),
	.dataf(!\always10~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always10),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~9 .extended_lut = "off";
defparam \always10~9 .lut_mask = 64'hAFAF008C00000000;
defparam \always10~9 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!comb),
	.datab(!burst_uncompress_busy),
	.datac(!mem_38_0),
	.datad(!source_addr_2),
	.datae(!mem_39_0),
	.dataf(!source_addr_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft0),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h4040000040FB00BB;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan15~0 (
	.dataa(!mem_124_0),
	.datab(!mem_122_0),
	.datac(!mem_123_0),
	.datad(!mem_90_0),
	.datae(!mem_91_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan15),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan15~0 .extended_lut = "off";
defparam \LessThan15~0 .lut_mask = 64'h80A0A8AA80A0A8AA;
defparam \LessThan15~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!comb),
	.datab(!burst_uncompress_busy),
	.datac(!mem_38_0),
	.datad(!source_addr_2),
	.datae(!mem_39_0),
	.dataf(!source_addr_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft01),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h04040000BF04BB00;
defparam \ShiftLeft0~1 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!comb),
	.datab(!burst_uncompress_busy),
	.datac(!mem_38_0),
	.datad(!source_addr_2),
	.datae(!mem_39_0),
	.dataf(!source_addr_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ShiftLeft02),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00BB40FB00004040;
defparam \ShiftLeft0~2 .shared_arith = "off";

cyclonev_lcell_comb \p1_ready~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!h2f_RREADY_0),
	.datac(!src0_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(p1_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \p1_ready~0 .extended_lut = "off";
defparam \p1_ready~0 .lut_mask = 64'h3535353535353535;
defparam \p1_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \always10~10 (
	.dataa(!src_payload),
	.datab(!always10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always101),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~10 .extended_lut = "off";
defparam \always10~10 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always10~10 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~0 (
	.dataa(!q_b_0),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_0_0),
	.datae(!data_reg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~0 .extended_lut = "off";
defparam \data_reg~0 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \always9~0 (
	.dataa(!h2f_BREADY_0),
	.datab(!h2f_RREADY_0),
	.datac(!out_valid),
	.datad(!src_payload),
	.datae(!always10),
	.dataf(!src0_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always9~0 .extended_lut = "off";
defparam \always9~0 .lut_mask = 64'h3030F0305050F050;
defparam \always9~0 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~1 (
	.dataa(!ShiftLeft0),
	.datab(!out_data_1),
	.datac(!data_reg_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~1 .extended_lut = "off";
defparam \data_reg~1 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~2 (
	.dataa(!q_b_2),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_2_0),
	.datae(!data_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~2 .extended_lut = "off";
defparam \data_reg~2 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~2 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~3 (
	.dataa(!q_b_3),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_3_0),
	.datae(!data_reg_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~3 .extended_lut = "off";
defparam \data_reg~3 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~4 (
	.dataa(!ShiftLeft0),
	.datab(!out_data_4),
	.datac(!data_reg_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~4 .extended_lut = "off";
defparam \data_reg~4 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~4 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~5 (
	.dataa(!q_b_5),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_5_0),
	.datae(!data_reg_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~5 .extended_lut = "off";
defparam \data_reg~5 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~5 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~6 (
	.dataa(!ShiftLeft0),
	.datab(!out_data_6),
	.datac(!data_reg_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~6 .extended_lut = "off";
defparam \data_reg~6 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~7 (
	.dataa(!q_b_7),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_7_0),
	.datae(!data_reg_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~7 .extended_lut = "off";
defparam \data_reg~7 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~7 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~8 (
	.dataa(!ShiftLeft0),
	.datab(!out_data_8),
	.datac(!data_reg_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~8 .extended_lut = "off";
defparam \data_reg~8 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~8 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~9 (
	.dataa(!q_b_9),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_9_0),
	.datae(!data_reg_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~9 .extended_lut = "off";
defparam \data_reg~9 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~9 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~10 (
	.dataa(!q_b_10),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_10_0),
	.datae(!data_reg_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~10 .extended_lut = "off";
defparam \data_reg~10 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~10 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~11 (
	.dataa(!q_b_11),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_11_0),
	.datae(!data_reg_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~11 .extended_lut = "off";
defparam \data_reg~11 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~11 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~12 (
	.dataa(!q_b_12),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_12_0),
	.datae(!data_reg_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~12 .extended_lut = "off";
defparam \data_reg~12 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~12 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~13 (
	.dataa(!ShiftLeft0),
	.datab(!out_data_13),
	.datac(!data_reg_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~13 .extended_lut = "off";
defparam \data_reg~13 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~13 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~14 (
	.dataa(!q_b_14),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_14_0),
	.datae(!data_reg_14),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~14 .extended_lut = "off";
defparam \data_reg~14 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~14 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~15 (
	.dataa(!q_b_15),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_15_0),
	.datae(!data_reg_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~15 .extended_lut = "off";
defparam \data_reg~15 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~15 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~16 (
	.dataa(!q_b_16),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_16_0),
	.datae(!data_reg_16),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~16 .extended_lut = "off";
defparam \data_reg~16 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~16 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~17 (
	.dataa(!ShiftLeft0),
	.datab(!out_data_17),
	.datac(!data_reg_17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~17 .extended_lut = "off";
defparam \data_reg~17 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~17 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~18 (
	.dataa(!q_b_18),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_18_0),
	.datae(!data_reg_18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~18 .extended_lut = "off";
defparam \data_reg~18 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~18 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~19 (
	.dataa(!q_b_19),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_19_0),
	.datae(!data_reg_19),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~19 .extended_lut = "off";
defparam \data_reg~19 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~19 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~20 (
	.dataa(!ShiftLeft0),
	.datab(!out_data_20),
	.datac(!data_reg_20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~20 .extended_lut = "off";
defparam \data_reg~20 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~20 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~21 (
	.dataa(!q_b_21),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_21_0),
	.datae(!data_reg_21),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~21 .extended_lut = "off";
defparam \data_reg~21 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~21 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~22 (
	.dataa(!ShiftLeft0),
	.datab(!out_data_22),
	.datac(!data_reg_22),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~22 .extended_lut = "off";
defparam \data_reg~22 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~22 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~23 (
	.dataa(!q_b_23),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_23_0),
	.datae(!data_reg_23),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~23 .extended_lut = "off";
defparam \data_reg~23 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~23 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~24 (
	.dataa(!ShiftLeft0),
	.datab(!out_data_24),
	.datac(!data_reg_24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~24 .extended_lut = "off";
defparam \data_reg~24 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~24 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~25 (
	.dataa(!q_b_25),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_25_0),
	.datae(!data_reg_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~25 .extended_lut = "off";
defparam \data_reg~25 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~25 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~26 (
	.dataa(!q_b_26),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_26_0),
	.datae(!data_reg_26),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~26 .extended_lut = "off";
defparam \data_reg~26 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~26 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~27 (
	.dataa(!q_b_27),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_27_0),
	.datae(!data_reg_27),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~27 .extended_lut = "off";
defparam \data_reg~27 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~27 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~28 (
	.dataa(!q_b_28),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_28_0),
	.datae(!data_reg_28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~28 .extended_lut = "off";
defparam \data_reg~28 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~28 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~29 (
	.dataa(!ShiftLeft0),
	.datab(!out_data_29),
	.datac(!data_reg_29),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~29 .extended_lut = "off";
defparam \data_reg~29 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~29 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~30 (
	.dataa(!q_b_30),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_30_0),
	.datae(!data_reg_30),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~30 .extended_lut = "off";
defparam \data_reg~30 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~30 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~31 (
	.dataa(!q_b_31),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_31_0),
	.datae(!data_reg_31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~31 .extended_lut = "off";
defparam \data_reg~31 .lut_mask = 64'h0131FFFF0131FFFF;
defparam \data_reg~31 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~32 (
	.dataa(!q_b_0),
	.datab(!always4),
	.datac(!mem_0_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_32),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~32 .extended_lut = "off";
defparam \data_reg~32 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~32 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~33 (
	.dataa(!out_data_1),
	.datab(!ShiftLeft01),
	.datac(!data_reg_33),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~33 .extended_lut = "off";
defparam \data_reg~33 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~33 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~34 (
	.dataa(!q_b_2),
	.datab(!always4),
	.datac(!mem_2_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_34),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~34 .extended_lut = "off";
defparam \data_reg~34 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~34 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~35 (
	.dataa(!q_b_3),
	.datab(!always4),
	.datac(!mem_3_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_35),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~35 .extended_lut = "off";
defparam \data_reg~35 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~35 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~36 (
	.dataa(!out_data_4),
	.datab(!ShiftLeft01),
	.datac(!data_reg_36),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~36 .extended_lut = "off";
defparam \data_reg~36 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~36 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~37 (
	.dataa(!q_b_5),
	.datab(!always4),
	.datac(!mem_5_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_37),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~37 .extended_lut = "off";
defparam \data_reg~37 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~37 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~38 (
	.dataa(!out_data_6),
	.datab(!ShiftLeft01),
	.datac(!data_reg_38),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~38 .extended_lut = "off";
defparam \data_reg~38 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~38 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~39 (
	.dataa(!q_b_7),
	.datab(!always4),
	.datac(!mem_7_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_39),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~39 .extended_lut = "off";
defparam \data_reg~39 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~39 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~40 (
	.dataa(!out_data_8),
	.datab(!ShiftLeft01),
	.datac(!data_reg_40),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~40 .extended_lut = "off";
defparam \data_reg~40 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~40 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~41 (
	.dataa(!q_b_9),
	.datab(!always4),
	.datac(!mem_9_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_41),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~41 .extended_lut = "off";
defparam \data_reg~41 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~41 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~42 (
	.dataa(!q_b_10),
	.datab(!always4),
	.datac(!mem_10_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_42),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~42 .extended_lut = "off";
defparam \data_reg~42 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~42 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~43 (
	.dataa(!q_b_11),
	.datab(!always4),
	.datac(!mem_11_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_43),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~43 .extended_lut = "off";
defparam \data_reg~43 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~43 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~44 (
	.dataa(!q_b_12),
	.datab(!always4),
	.datac(!mem_12_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_44),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~44 .extended_lut = "off";
defparam \data_reg~44 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~44 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~45 (
	.dataa(!out_data_13),
	.datab(!ShiftLeft01),
	.datac(!data_reg_45),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~45 .extended_lut = "off";
defparam \data_reg~45 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~45 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~46 (
	.dataa(!q_b_14),
	.datab(!always4),
	.datac(!mem_14_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_46),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~46 .extended_lut = "off";
defparam \data_reg~46 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~46 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~47 (
	.dataa(!q_b_15),
	.datab(!always4),
	.datac(!mem_15_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_47),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~47 .extended_lut = "off";
defparam \data_reg~47 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~47 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~48 (
	.dataa(!q_b_16),
	.datab(!always4),
	.datac(!mem_16_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_48),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~48 .extended_lut = "off";
defparam \data_reg~48 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~48 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~49 (
	.dataa(!out_data_17),
	.datab(!ShiftLeft01),
	.datac(!data_reg_49),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~49 .extended_lut = "off";
defparam \data_reg~49 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~49 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~50 (
	.dataa(!q_b_18),
	.datab(!always4),
	.datac(!mem_18_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_50),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~50 .extended_lut = "off";
defparam \data_reg~50 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~50 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~51 (
	.dataa(!q_b_19),
	.datab(!always4),
	.datac(!mem_19_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_51),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~51 .extended_lut = "off";
defparam \data_reg~51 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~51 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~52 (
	.dataa(!out_data_20),
	.datab(!ShiftLeft01),
	.datac(!data_reg_52),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~52 .extended_lut = "off";
defparam \data_reg~52 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~52 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~53 (
	.dataa(!q_b_21),
	.datab(!always4),
	.datac(!mem_21_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_53),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~53 .extended_lut = "off";
defparam \data_reg~53 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~53 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~54 (
	.dataa(!out_data_22),
	.datab(!ShiftLeft01),
	.datac(!data_reg_54),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~54 .extended_lut = "off";
defparam \data_reg~54 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~54 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~55 (
	.dataa(!q_b_23),
	.datab(!always4),
	.datac(!mem_23_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_55),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~55 .extended_lut = "off";
defparam \data_reg~55 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~55 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~56 (
	.dataa(!out_data_24),
	.datab(!ShiftLeft01),
	.datac(!data_reg_56),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~56 .extended_lut = "off";
defparam \data_reg~56 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~56 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~57 (
	.dataa(!q_b_25),
	.datab(!always4),
	.datac(!mem_25_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_57),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~57 .extended_lut = "off";
defparam \data_reg~57 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~57 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~58 (
	.dataa(!q_b_26),
	.datab(!always4),
	.datac(!mem_26_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_58),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~58 .extended_lut = "off";
defparam \data_reg~58 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~58 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~59 (
	.dataa(!q_b_27),
	.datab(!always4),
	.datac(!mem_27_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_59),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~59 .extended_lut = "off";
defparam \data_reg~59 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~59 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~60 (
	.dataa(!q_b_28),
	.datab(!always4),
	.datac(!mem_28_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_60),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~60 .extended_lut = "off";
defparam \data_reg~60 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~60 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~61 (
	.dataa(!out_data_29),
	.datab(!ShiftLeft01),
	.datac(!data_reg_61),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~61 .extended_lut = "off";
defparam \data_reg~61 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~61 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~62 (
	.dataa(!q_b_30),
	.datab(!always4),
	.datac(!mem_30_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_62),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~62 .extended_lut = "off";
defparam \data_reg~62 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~62 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~63 (
	.dataa(!q_b_31),
	.datab(!always4),
	.datac(!mem_31_0),
	.datad(!ShiftLeft01),
	.datae(!data_reg_63),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~63 .extended_lut = "off";
defparam \data_reg~63 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~63 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~64 (
	.dataa(!q_b_0),
	.datab(!always4),
	.datac(!mem_0_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_64),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~64 .extended_lut = "off";
defparam \data_reg~64 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~64 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~65 (
	.dataa(!out_data_1),
	.datab(!ShiftLeft02),
	.datac(!data_reg_65),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~65 .extended_lut = "off";
defparam \data_reg~65 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~65 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~66 (
	.dataa(!q_b_2),
	.datab(!always4),
	.datac(!mem_2_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_66),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~66 .extended_lut = "off";
defparam \data_reg~66 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~66 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~67 (
	.dataa(!q_b_3),
	.datab(!always4),
	.datac(!mem_3_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_67),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~67 .extended_lut = "off";
defparam \data_reg~67 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~67 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~68 (
	.dataa(!out_data_4),
	.datab(!ShiftLeft02),
	.datac(!data_reg_68),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~68 .extended_lut = "off";
defparam \data_reg~68 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~68 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~69 (
	.dataa(!q_b_5),
	.datab(!always4),
	.datac(!mem_5_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_69),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~69 .extended_lut = "off";
defparam \data_reg~69 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~69 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~70 (
	.dataa(!out_data_6),
	.datab(!ShiftLeft02),
	.datac(!data_reg_70),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~70 .extended_lut = "off";
defparam \data_reg~70 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~70 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~71 (
	.dataa(!q_b_7),
	.datab(!always4),
	.datac(!mem_7_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_71),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~71_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~71 .extended_lut = "off";
defparam \data_reg~71 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~71 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~72 (
	.dataa(!out_data_8),
	.datab(!ShiftLeft02),
	.datac(!data_reg_72),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~72 .extended_lut = "off";
defparam \data_reg~72 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~72 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~73 (
	.dataa(!q_b_9),
	.datab(!always4),
	.datac(!mem_9_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_73),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~73 .extended_lut = "off";
defparam \data_reg~73 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~73 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~74 (
	.dataa(!q_b_10),
	.datab(!always4),
	.datac(!mem_10_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_74),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~74_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~74 .extended_lut = "off";
defparam \data_reg~74 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~74 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~75 (
	.dataa(!q_b_11),
	.datab(!always4),
	.datac(!mem_11_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_75),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~75_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~75 .extended_lut = "off";
defparam \data_reg~75 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~75 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~76 (
	.dataa(!q_b_12),
	.datab(!always4),
	.datac(!mem_12_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_76),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~76_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~76 .extended_lut = "off";
defparam \data_reg~76 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~76 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~77 (
	.dataa(!out_data_13),
	.datab(!ShiftLeft02),
	.datac(!data_reg_77),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~77_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~77 .extended_lut = "off";
defparam \data_reg~77 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~77 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~78 (
	.dataa(!q_b_14),
	.datab(!always4),
	.datac(!mem_14_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_78),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~78_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~78 .extended_lut = "off";
defparam \data_reg~78 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~78 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~79 (
	.dataa(!q_b_15),
	.datab(!always4),
	.datac(!mem_15_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_79),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~79_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~79 .extended_lut = "off";
defparam \data_reg~79 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~79 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~80 (
	.dataa(!q_b_16),
	.datab(!always4),
	.datac(!mem_16_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_80),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~80_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~80 .extended_lut = "off";
defparam \data_reg~80 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~80 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~81 (
	.dataa(!out_data_17),
	.datab(!ShiftLeft02),
	.datac(!data_reg_81),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~81_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~81 .extended_lut = "off";
defparam \data_reg~81 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~81 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~82 (
	.dataa(!q_b_18),
	.datab(!always4),
	.datac(!mem_18_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_82),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~82_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~82 .extended_lut = "off";
defparam \data_reg~82 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~82 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~83 (
	.dataa(!q_b_19),
	.datab(!always4),
	.datac(!mem_19_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_83),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~83_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~83 .extended_lut = "off";
defparam \data_reg~83 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~83 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~84 (
	.dataa(!out_data_20),
	.datab(!ShiftLeft02),
	.datac(!data_reg_84),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~84_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~84 .extended_lut = "off";
defparam \data_reg~84 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~84 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~85 (
	.dataa(!q_b_21),
	.datab(!always4),
	.datac(!mem_21_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_85),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~85_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~85 .extended_lut = "off";
defparam \data_reg~85 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~85 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~86 (
	.dataa(!out_data_22),
	.datab(!ShiftLeft02),
	.datac(!data_reg_86),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~86_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~86 .extended_lut = "off";
defparam \data_reg~86 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~86 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~87 (
	.dataa(!q_b_23),
	.datab(!always4),
	.datac(!mem_23_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_87),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~87_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~87 .extended_lut = "off";
defparam \data_reg~87 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~87 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~88 (
	.dataa(!out_data_24),
	.datab(!ShiftLeft02),
	.datac(!data_reg_88),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~88_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~88 .extended_lut = "off";
defparam \data_reg~88 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~88 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~89 (
	.dataa(!q_b_25),
	.datab(!always4),
	.datac(!mem_25_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_89),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~89_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~89 .extended_lut = "off";
defparam \data_reg~89 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~89 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~90 (
	.dataa(!q_b_26),
	.datab(!always4),
	.datac(!mem_26_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_90),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~90_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~90 .extended_lut = "off";
defparam \data_reg~90 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~90 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~91 (
	.dataa(!q_b_27),
	.datab(!always4),
	.datac(!mem_27_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_91),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~91_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~91 .extended_lut = "off";
defparam \data_reg~91 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~91 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~92 (
	.dataa(!q_b_28),
	.datab(!always4),
	.datac(!mem_28_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_92),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~92_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~92 .extended_lut = "off";
defparam \data_reg~92 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~92 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~93 (
	.dataa(!out_data_29),
	.datab(!ShiftLeft02),
	.datac(!data_reg_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~93_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~93 .extended_lut = "off";
defparam \data_reg~93 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \data_reg~93 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~94 (
	.dataa(!q_b_30),
	.datab(!always4),
	.datac(!mem_30_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_94),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~94_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~94 .extended_lut = "off";
defparam \data_reg~94 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~94 .shared_arith = "off";

cyclonev_lcell_comb \data_reg~95 (
	.dataa(!q_b_31),
	.datab(!always4),
	.datac(!mem_31_0),
	.datad(!ShiftLeft02),
	.datae(!data_reg_95),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_reg~95_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_reg~95 .extended_lut = "off";
defparam \data_reg~95 .lut_mask = 64'h001DFFFF001DFFFF;
defparam \data_reg~95 .shared_arith = "off";

cyclonev_lcell_comb \always10~0 (
	.dataa(!mem_123_0),
	.datab(!mem_91_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~0 .extended_lut = "off";
defparam \always10~0 .lut_mask = 64'h4444444444444444;
defparam \always10~0 .shared_arith = "off";

cyclonev_lcell_comb \always10~1 (
	.dataa(!comb),
	.datab(!mem_122_0),
	.datac(!burst_uncompress_busy),
	.datad(!mem_38_0),
	.datae(!source_addr_2),
	.dataf(!\always10~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~1 .extended_lut = "off";
defparam \always10~1 .lut_mask = 64'hEFFFCCDC00000000;
defparam \always10~1 .shared_arith = "off";

cyclonev_lcell_comb \ShiftRight0~0 (
	.dataa(!mem_122_0),
	.datab(!mem_123_0),
	.datac(!mem_124_0),
	.datad(!mem_90_0),
	.datae(!mem_91_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftRight0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftRight0~0 .extended_lut = "off";
defparam \ShiftRight0~0 .lut_mask = 64'h0804020108040201;
defparam \ShiftRight0~0 .shared_arith = "off";

cyclonev_lcell_comb \always10~2 (
	.dataa(!mem_122_0),
	.datab(!mem_123_0),
	.datac(!mem_90_0),
	.datad(!mem_91_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~2 .extended_lut = "off";
defparam \always10~2 .lut_mask = 64'h0008000800080008;
defparam \always10~2 .shared_arith = "off";

cyclonev_lcell_comb \always10~3 (
	.dataa(!comb),
	.datab(!\ShiftRight0~0_combout ),
	.datac(!burst_uncompress_busy),
	.datad(!mem_39_0),
	.datae(!source_addr_3),
	.dataf(!\always10~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~3 .extended_lut = "off";
defparam \always10~3 .lut_mask = 64'h5000FFAF10003323;
defparam \always10~3 .shared_arith = "off";

cyclonev_lcell_comb \always10~4 (
	.dataa(!mem_123_0),
	.datab(!mem_91_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~4 .extended_lut = "off";
defparam \always10~4 .lut_mask = 64'h2222222222222222;
defparam \always10~4 .shared_arith = "off";

cyclonev_lcell_comb \always10~5 (
	.dataa(!mem_122_0),
	.datab(!mem_90_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~5 .extended_lut = "off";
defparam \always10~5 .lut_mask = 64'h2222222222222222;
defparam \always10~5 .shared_arith = "off";

cyclonev_lcell_comb \always10~6 (
	.dataa(!comb),
	.datab(!burst_uncompress_busy),
	.datac(!mem_38_0),
	.datad(!source_addr_2),
	.datae(!\always10~4_combout ),
	.dataf(!\always10~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~6 .extended_lut = "off";
defparam \always10~6 .lut_mask = 64'hFFFF000040FB0000;
defparam \always10~6 .shared_arith = "off";

cyclonev_lcell_comb \always10~7 (
	.dataa(!mem_124_0),
	.datab(!\ShiftRight0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~7 .extended_lut = "off";
defparam \always10~7 .lut_mask = 64'h8888888888888888;
defparam \always10~7 .shared_arith = "off";

cyclonev_lcell_comb \always10~8 (
	.dataa(!mem_122_0),
	.datab(!mem_123_0),
	.datac(!mem_90_0),
	.datad(!mem_91_0),
	.datae(!\ShiftRight0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~8 .extended_lut = "off";
defparam \always10~8 .lut_mask = 64'h8421000084210000;
defparam \always10~8 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_cmd_demux (
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	in_ready_hold,
	saved_grant_0,
	in_ready,
	nxt_in_ready,
	nxt_in_ready1,
	Equal0,
	Equal01,
	Equal02,
	sink_ready,
	nxt_in_ready2,
	load_next_out_cmd,
	Equal03,
	saved_grant_01,
	count_1,
	count_0,
	sink_ready1,
	last_channel_0,
	has_pending_responses,
	last_cycle,
	last_channel_1,
	src1_valid,
	src0_valid,
	sink_ready2,
	src0_valid1,
	sink_ready3)/* synthesis synthesis_greybox=0 */;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	in_ready_hold;
input 	saved_grant_0;
input 	in_ready;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	Equal0;
input 	Equal01;
input 	Equal02;
output 	sink_ready;
input 	nxt_in_ready2;
input 	load_next_out_cmd;
input 	Equal03;
input 	saved_grant_01;
input 	count_1;
input 	count_0;
output 	sink_ready1;
input 	last_channel_0;
input 	has_pending_responses;
input 	last_cycle;
input 	last_channel_1;
output 	src1_valid;
output 	src0_valid;
output 	sink_ready2;
output 	src0_valid1;
output 	sink_ready3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~1_combout ;


cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!saved_grant_0),
	.datab(!Equal0),
	.datac(!Equal01),
	.datad(!Equal02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h5554555455545554;
defparam \sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~2 (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready2),
	.datac(!load_next_out_cmd),
	.datad(!Equal0),
	.datae(!Equal03),
	.dataf(!\sink_ready~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~2 .extended_lut = "off";
defparam \sink_ready~2 .lut_mask = 64'h000000000000001D;
defparam \sink_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!has_pending_responses),
	.datab(!last_cycle),
	.datac(!last_channel_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h2323232323232323;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!last_channel_0),
	.datab(!has_pending_responses),
	.datac(!last_cycle),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'h0D0D0D0D0D0D0D0D;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~3 (
	.dataa(!in_ready),
	.datab(!nxt_in_ready),
	.datac(!nxt_in_ready1),
	.datad(!sink_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~3 .extended_lut = "off";
defparam \sink_ready~3 .lut_mask = 64'h00A200A200A200A2;
defparam \sink_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~1 (
	.dataa(!Equal0),
	.datab(!Equal01),
	.datac(!Equal02),
	.datad(!src0_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~1 .extended_lut = "off";
defparam \src0_valid~1 .lut_mask = 64'h0001000100010001;
defparam \src0_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~4 (
	.dataa(!Equal0),
	.datab(!Equal01),
	.datac(!Equal02),
	.datad(!\sink_ready~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready3),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~4 .extended_lut = "off";
defparam \sink_ready~4 .lut_mask = 64'h0001000100010001;
defparam \sink_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~1 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!h2f_AWSIZE_1),
	.datac(!h2f_AWSIZE_2),
	.datad(!saved_grant_01),
	.datae(!count_1),
	.dataf(!count_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~1 .extended_lut = "off";
defparam \sink_ready~1 .lut_mask = 64'h00E000E000FF00E0;
defparam \sink_ready~1 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_cmd_mux (
	h2f_AWVALID_0,
	h2f_WLAST_0,
	h2f_WVALID_0,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	outclk_wire_0,
	in_ready_hold,
	Equal0,
	Equal01,
	Equal02,
	nxt_in_ready,
	load_next_out_cmd,
	Equal03,
	saved_grant_0,
	sink_ready,
	last_channel_0,
	has_pending_responses,
	last_cycle,
	last_cycle1,
	r_sync_rst,
	src0_valid,
	src_payload,
	src_payload1,
	src_payload2,
	Selector7,
	nxt_in_ready1,
	nxt_in_ready2,
	src0_valid1,
	sink_ready1,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15)/* synthesis synthesis_greybox=0 */;
input 	h2f_AWVALID_0;
input 	h2f_WLAST_0;
input 	h2f_WVALID_0;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	outclk_wire_0;
input 	in_ready_hold;
input 	Equal0;
input 	Equal01;
input 	Equal02;
input 	nxt_in_ready;
input 	load_next_out_cmd;
input 	Equal03;
output 	saved_grant_0;
input 	sink_ready;
input 	last_channel_0;
input 	has_pending_responses;
output 	last_cycle;
output 	last_cycle1;
input 	r_sync_rst;
input 	src0_valid;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
input 	Selector7;
input 	nxt_in_ready1;
input 	nxt_in_ready2;
input 	src0_valid1;
input 	sink_ready1;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \last_cycle~2_combout ;
wire \update_grant~1_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \saved_grant[0]~0_combout ;


Computer_System_altera_merlin_arbitrator_1 arb(
	.clk(outclk_wire_0),
	.Equal0(Equal0),
	.Equal01(Equal03),
	.reset(r_sync_rst),
	.src0_valid(src0_valid),
	.update_grant(\update_grant~0_combout ),
	.last_cycle(\last_cycle~2_combout ),
	.grant_0(\arb|grant[0]~0_combout ),
	.nxt_in_ready(nxt_in_ready1),
	.nxt_in_ready1(nxt_in_ready2),
	.src0_valid1(src0_valid1),
	.sink_ready(sink_ready1));

dffeas \saved_grant[0] (
	.clk(outclk_wire_0),
	.d(\saved_grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \last_cycle~0 (
	.dataa(!h2f_AWVALID_0),
	.datab(!h2f_WLAST_0),
	.datac(!h2f_WVALID_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_cycle),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_cycle~0 .extended_lut = "off";
defparam \last_cycle~0 .lut_mask = 64'h0101010101010101;
defparam \last_cycle~0 .shared_arith = "off";

cyclonev_lcell_comb \last_cycle~1 (
	.dataa(!h2f_AWVALID_0),
	.datab(!h2f_WVALID_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_cycle1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_cycle~1 .extended_lut = "off";
defparam \last_cycle~1 .lut_mask = 64'h1111111111111111;
defparam \last_cycle~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_AWSIZE_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_AWSIZE_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_AWSIZE_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!h2f_AWID_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h1111111111111111;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!h2f_AWID_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1111111111111111;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!h2f_AWID_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h1111111111111111;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!h2f_AWID_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h1111111111111111;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!h2f_AWID_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h1111111111111111;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!h2f_AWID_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h1111111111111111;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!h2f_AWID_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h1111111111111111;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!h2f_AWID_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h1111111111111111;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!h2f_AWID_8),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h1111111111111111;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!h2f_AWID_9),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h1111111111111111;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!h2f_AWID_10),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h1111111111111111;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!h2f_AWID_11),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h1111111111111111;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!Selector7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h4444444444444444;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \last_cycle~2 (
	.dataa(!last_channel_0),
	.datab(!has_pending_responses),
	.datac(!last_cycle),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_cycle~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_cycle~2 .extended_lut = "off";
defparam \last_cycle~2 .lut_mask = 64'h0D0D0D0D0D0D0D0D;
defparam \last_cycle~2 .shared_arith = "off";

cyclonev_lcell_comb \update_grant~1 (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready),
	.datac(!load_next_out_cmd),
	.datad(!sink_ready1),
	.datae(!\update_grant~0_combout ),
	.dataf(!\last_cycle~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~1 .extended_lut = "off";
defparam \update_grant~1 .lut_mask = 64'hFFFF0000FFE20000;
defparam \update_grant~1 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(outclk_wire_0),
	.d(\update_grant~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!Equal0),
	.datac(!Equal01),
	.datad(!Equal02),
	.datae(!\packet_in_progress~q ),
	.dataf(!src0_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFFFF0000FFFE0000;
defparam \update_grant~0 .shared_arith = "off";

cyclonev_lcell_comb \saved_grant[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!sink_ready),
	.datac(!\update_grant~0_combout ),
	.datad(!\last_cycle~2_combout ),
	.datae(!\arb|grant[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[0]~0 .extended_lut = "off";
defparam \saved_grant[0]~0 .lut_mask = 64'h50405F7F50405F7F;
defparam \saved_grant[0]~0 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_cmd_mux_1 (
	h2f_WLAST_0,
	h2f_ARADDR_0,
	h2f_ARADDR_2,
	h2f_ARADDR_4,
	h2f_ARADDR_5,
	h2f_ARADDR_6,
	h2f_ARADDR_7,
	h2f_ARADDR_8,
	h2f_ARADDR_9,
	h2f_ARBURST_0,
	h2f_ARBURST_1,
	h2f_ARID_0,
	h2f_ARID_1,
	h2f_ARID_2,
	h2f_ARID_3,
	h2f_ARID_4,
	h2f_ARID_5,
	h2f_ARID_6,
	h2f_ARID_7,
	h2f_ARID_8,
	h2f_ARID_9,
	h2f_ARID_10,
	h2f_ARID_11,
	h2f_ARLEN_0,
	h2f_ARLEN_1,
	h2f_ARLEN_2,
	h2f_ARLEN_3,
	h2f_ARSIZE_0,
	h2f_ARSIZE_1,
	h2f_ARSIZE_2,
	h2f_AWADDR_0,
	h2f_AWBURST_0,
	h2f_AWBURST_1,
	h2f_AWID_0,
	h2f_AWID_1,
	h2f_AWID_2,
	h2f_AWID_3,
	h2f_AWID_4,
	h2f_AWID_5,
	h2f_AWID_6,
	h2f_AWID_7,
	h2f_AWID_8,
	h2f_AWID_9,
	h2f_AWID_10,
	h2f_AWID_11,
	h2f_AWLEN_0,
	h2f_AWLEN_1,
	h2f_AWLEN_2,
	h2f_AWSIZE_0,
	h2f_AWSIZE_1,
	h2f_AWSIZE_2,
	h2f_WSTRB_0,
	h2f_WSTRB_1,
	h2f_WSTRB_2,
	h2f_WSTRB_3,
	h2f_WSTRB_4,
	h2f_WSTRB_5,
	h2f_WSTRB_6,
	h2f_WSTRB_7,
	h2f_WSTRB_8,
	h2f_WSTRB_9,
	h2f_WSTRB_10,
	h2f_WSTRB_11,
	h2f_WSTRB_12,
	h2f_WSTRB_13,
	h2f_WSTRB_14,
	h2f_WSTRB_15,
	outclk_wire_0,
	Add4,
	Add5,
	Add41,
	Add51,
	Add42,
	Add52,
	Add43,
	Add53,
	Add44,
	Add54,
	Add55,
	Add45,
	Add56,
	Add46,
	Add47,
	Add57,
	Add48,
	Add58,
	src_data_185,
	saved_grant_1,
	saved_grant_0,
	src_data_198,
	src_data_199,
	src_data_200,
	in_ready,
	nxt_in_ready,
	nxt_in_ready1,
	sink1_ready1,
	nxt_in_ready2,
	sop_enable,
	Equal0,
	Equal01,
	Equal02,
	r_sync_rst,
	Equal03,
	cmd_src_valid_1,
	src1_valid,
	WideOr11,
	src_payload_0,
	LessThan11,
	src_payload,
	Add3,
	log2ceil,
	src_data_190,
	LessThan10,
	src_payload1,
	Add31,
	src_data_189,
	address_burst_0,
	src_data_144,
	src_data_130,
	src_data_134,
	src_data_138,
	src_data_142,
	out_data_2,
	src_data_146,
	src_data_128,
	src_data_132,
	src_data_136,
	src_data_140,
	src_data_129,
	src_data_133,
	src_data_137,
	src_data_141,
	src_data_131,
	src_data_135,
	src_data_139,
	src_data_143,
	burst_bytecount_4,
	src_data_184,
	burst_bytecount_6,
	src_payload2,
	src_payload3,
	burst_bytecount_5,
	src_payload4,
	src_payload5,
	burst_bytecount_7,
	Add0,
	Add2,
	src_data_187,
	Add01,
	Add21,
	src_data_186,
	Add22,
	write_cp_data_188,
	src_payload6,
	src_data_188,
	src_payload7,
	src_valid,
	Add1,
	out_data_9,
	LessThan16,
	out_data_8,
	LessThan12,
	Selector26,
	LessThan14,
	LessThan15,
	src_payload8,
	src_data_191,
	src_payload9,
	src_data_192,
	src_data_193,
	src_data_1931,
	src_payload10,
	src_data_194,
	src_data_1941,
	src_payload11,
	src_data_195,
	src_data_1951,
	src_payload12,
	src_data_196,
	Add32,
	src_data_1961,
	src_payload13,
	src_data_197,
	src_data_1971,
	src_data_152,
	src_payload14,
	src_payload15,
	Selector7,
	src_data_1901,
	Selector8,
	src_data_1891,
	src_data_209,
	src_data_210,
	src_data_211,
	src_data_212,
	src_data_213,
	src_data_214,
	src_data_215,
	src_data_216,
	src_data_217,
	src_data_218,
	src_data_219,
	src_data_220,
	Selector6,
	src_data_1911,
	Selector5,
	src_data_1921,
	src_data_1932,
	src_data_1942,
	src_data_1952,
	src_data_1962,
	src_data_1972)/* synthesis synthesis_greybox=0 */;
input 	h2f_WLAST_0;
input 	h2f_ARADDR_0;
input 	h2f_ARADDR_2;
input 	h2f_ARADDR_4;
input 	h2f_ARADDR_5;
input 	h2f_ARADDR_6;
input 	h2f_ARADDR_7;
input 	h2f_ARADDR_8;
input 	h2f_ARADDR_9;
input 	h2f_ARBURST_0;
input 	h2f_ARBURST_1;
input 	h2f_ARID_0;
input 	h2f_ARID_1;
input 	h2f_ARID_2;
input 	h2f_ARID_3;
input 	h2f_ARID_4;
input 	h2f_ARID_5;
input 	h2f_ARID_6;
input 	h2f_ARID_7;
input 	h2f_ARID_8;
input 	h2f_ARID_9;
input 	h2f_ARID_10;
input 	h2f_ARID_11;
input 	h2f_ARLEN_0;
input 	h2f_ARLEN_1;
input 	h2f_ARLEN_2;
input 	h2f_ARLEN_3;
input 	h2f_ARSIZE_0;
input 	h2f_ARSIZE_1;
input 	h2f_ARSIZE_2;
input 	h2f_AWADDR_0;
input 	h2f_AWBURST_0;
input 	h2f_AWBURST_1;
input 	h2f_AWID_0;
input 	h2f_AWID_1;
input 	h2f_AWID_2;
input 	h2f_AWID_3;
input 	h2f_AWID_4;
input 	h2f_AWID_5;
input 	h2f_AWID_6;
input 	h2f_AWID_7;
input 	h2f_AWID_8;
input 	h2f_AWID_9;
input 	h2f_AWID_10;
input 	h2f_AWID_11;
input 	h2f_AWLEN_0;
input 	h2f_AWLEN_1;
input 	h2f_AWLEN_2;
input 	h2f_AWSIZE_0;
input 	h2f_AWSIZE_1;
input 	h2f_AWSIZE_2;
input 	h2f_WSTRB_0;
input 	h2f_WSTRB_1;
input 	h2f_WSTRB_2;
input 	h2f_WSTRB_3;
input 	h2f_WSTRB_4;
input 	h2f_WSTRB_5;
input 	h2f_WSTRB_6;
input 	h2f_WSTRB_7;
input 	h2f_WSTRB_8;
input 	h2f_WSTRB_9;
input 	h2f_WSTRB_10;
input 	h2f_WSTRB_11;
input 	h2f_WSTRB_12;
input 	h2f_WSTRB_13;
input 	h2f_WSTRB_14;
input 	h2f_WSTRB_15;
input 	outclk_wire_0;
input 	Add4;
input 	Add5;
input 	Add41;
input 	Add51;
input 	Add42;
input 	Add52;
input 	Add43;
input 	Add53;
input 	Add44;
input 	Add54;
input 	Add55;
input 	Add45;
input 	Add56;
input 	Add46;
input 	Add47;
input 	Add57;
input 	Add48;
input 	Add58;
output 	src_data_185;
output 	saved_grant_1;
output 	saved_grant_0;
output 	src_data_198;
output 	src_data_199;
output 	src_data_200;
input 	in_ready;
input 	nxt_in_ready;
input 	nxt_in_ready1;
output 	sink1_ready1;
input 	nxt_in_ready2;
input 	sop_enable;
input 	Equal0;
input 	Equal01;
input 	Equal02;
input 	r_sync_rst;
input 	Equal03;
input 	cmd_src_valid_1;
input 	src1_valid;
output 	WideOr11;
output 	src_payload_0;
input 	LessThan11;
output 	src_payload;
input 	Add3;
input 	log2ceil;
output 	src_data_190;
input 	LessThan10;
output 	src_payload1;
input 	Add31;
output 	src_data_189;
input 	address_burst_0;
output 	src_data_144;
output 	src_data_130;
output 	src_data_134;
output 	src_data_138;
output 	src_data_142;
input 	out_data_2;
output 	src_data_146;
output 	src_data_128;
output 	src_data_132;
output 	src_data_136;
output 	src_data_140;
output 	src_data_129;
output 	src_data_133;
output 	src_data_137;
output 	src_data_141;
output 	src_data_131;
output 	src_data_135;
output 	src_data_139;
output 	src_data_143;
input 	burst_bytecount_4;
output 	src_data_184;
input 	burst_bytecount_6;
output 	src_payload2;
output 	src_payload3;
input 	burst_bytecount_5;
output 	src_payload4;
output 	src_payload5;
input 	burst_bytecount_7;
input 	Add0;
input 	Add2;
output 	src_data_187;
input 	Add01;
input 	Add21;
output 	src_data_186;
input 	Add22;
input 	write_cp_data_188;
output 	src_payload6;
output 	src_data_188;
output 	src_payload7;
output 	src_valid;
input 	Add1;
input 	out_data_9;
input 	LessThan16;
input 	out_data_8;
input 	LessThan12;
input 	Selector26;
input 	LessThan14;
input 	LessThan15;
output 	src_payload8;
output 	src_data_191;
output 	src_payload9;
output 	src_data_192;
output 	src_data_193;
output 	src_data_1931;
output 	src_payload10;
output 	src_data_194;
output 	src_data_1941;
output 	src_payload11;
output 	src_data_195;
output 	src_data_1951;
output 	src_payload12;
output 	src_data_196;
input 	Add32;
output 	src_data_1961;
output 	src_payload13;
output 	src_data_197;
output 	src_data_1971;
output 	src_data_152;
output 	src_payload14;
output 	src_payload15;
input 	Selector7;
output 	src_data_1901;
input 	Selector8;
output 	src_data_1891;
output 	src_data_209;
output 	src_data_210;
output 	src_data_211;
output 	src_data_212;
output 	src_data_213;
output 	src_data_214;
output 	src_data_215;
output 	src_data_216;
output 	src_data_217;
output 	src_data_218;
output 	src_data_219;
output 	src_data_220;
input 	Selector6;
output 	src_data_1911;
input 	Selector5;
output 	src_data_1921;
output 	src_data_1932;
output 	src_data_1942;
output 	src_data_1952;
output 	src_data_1962;
output 	src_data_1972;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \src_valid~0_combout ;
wire \src_data[190]~0_combout ;
wire \src_data[189]~2_combout ;
wire \src_data[189]~3_combout ;
wire \src_data[191]~5_combout ;
wire \src_data[193]~9_combout ;
wire \src_data[194]~11_combout ;
wire \src_data[195]~14_combout ;
wire \src_data[190]~21_combout ;
wire \src_data[189]~23_combout ;
wire \src_data[191]~25_combout ;
wire \src_data[192]~27_combout ;
wire \src_data[193]~29_combout ;
wire \src_data[193]~30_combout ;
wire \src_data[194]~32_combout ;
wire \src_data[194]~33_combout ;
wire \src_data[195]~35_combout ;
wire \src_data[195]~36_combout ;
wire \src_data[196]~38_combout ;
wire \src_data[196]~39_combout ;
wire \src_data[197]~41_combout ;


Computer_System_altera_merlin_arbitrator arb(
	.clk(outclk_wire_0),
	.in_ready(in_ready),
	.nxt_in_ready(nxt_in_ready2),
	.Equal0(Equal0),
	.Equal01(Equal01),
	.Equal02(Equal02),
	.reset(r_sync_rst),
	.Equal03(Equal03),
	.cmd_src_valid_1(cmd_src_valid_1),
	.src1_valid(src1_valid),
	.grant_1(\arb|grant[1]~0_combout ),
	.WideOr1(WideOr11),
	.src_payload_0(src_payload_0),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ));

cyclonev_lcell_comb \src_data[185]~43 (
	.dataa(!h2f_AWLEN_0),
	.datab(!Add22),
	.datac(!burst_bytecount_5),
	.datad(!saved_grant_0),
	.datae(!sop_enable),
	.dataf(!saved_grant_1),
	.datag(!h2f_AWLEN_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_185),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[185]~43 .extended_lut = "on";
defparam \src_data[185]~43 .lut_mask = 64'h005A000F337B333F;
defparam \src_data[185]~43 .shared_arith = "off";

dffeas \saved_grant[1] (
	.clk(outclk_wire_0),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(outclk_wire_0),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_data[198] (
	.dataa(!h2f_ARSIZE_0),
	.datab(!h2f_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_198),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[198] .extended_lut = "off";
defparam \src_data[198] .lut_mask = 64'h0537053705370537;
defparam \src_data[198] .shared_arith = "off";

cyclonev_lcell_comb \src_data[199] (
	.dataa(!h2f_ARSIZE_1),
	.datab(!h2f_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_199),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[199] .extended_lut = "off";
defparam \src_data[199] .lut_mask = 64'h0537053705370537;
defparam \src_data[199] .shared_arith = "off";

cyclonev_lcell_comb \src_data[200] (
	.dataa(!h2f_ARSIZE_2),
	.datab(!h2f_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_200),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[200] .extended_lut = "off";
defparam \src_data[200] .lut_mask = 64'h0537053705370537;
defparam \src_data[200] .shared_arith = "off";

cyclonev_lcell_comb sink1_ready(
	.dataa(!saved_grant_1),
	.datab(!in_ready),
	.datac(!nxt_in_ready),
	.datad(!nxt_in_ready1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink1_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam sink1_ready.extended_lut = "off";
defparam sink1_ready.lut_mask = 64'h4404440444044404;
defparam sink1_ready.shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!saved_grant_0),
	.datab(!Equal0),
	.datac(!Equal01),
	.datad(!Equal02),
	.datae(!src1_valid),
	.dataf(!\src_valid~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h00005554FFFFFFFF;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!saved_grant_0),
	.datad(!LessThan11),
	.datae(!Add4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h07050F0D07050F0D;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[190]~1 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!saved_grant_1),
	.datad(!Add5),
	.datae(!\src_data[190]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_190),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[190]~1 .extended_lut = "off";
defparam \src_data[190]~1 .lut_mask = 64'h070F050D070F050D;
defparam \src_data[190]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!saved_grant_0),
	.datad(!LessThan10),
	.datae(!Add41),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h07050F0D07050F0D;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[189]~4 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!saved_grant_1),
	.datad(!\src_data[189]~2_combout ),
	.datae(!Add51),
	.dataf(!\src_data[189]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_189),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[189]~4 .extended_lut = "off";
defparam \src_data[189]~4 .lut_mask = 64'h07070F0F07050F0D;
defparam \src_data[189]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[144] (
	.dataa(!h2f_ARADDR_0),
	.datab(!h2f_AWADDR_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(!sop_enable),
	.dataf(!address_burst_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_144),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[144] .extended_lut = "off";
defparam \src_data[144] .lut_mask = 64'h05370505053705FF;
defparam \src_data[144] .shared_arith = "off";

cyclonev_lcell_comb \src_data[130] (
	.dataa(!h2f_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_130),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[130] .extended_lut = "off";
defparam \src_data[130] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[130] .shared_arith = "off";

cyclonev_lcell_comb \src_data[134] (
	.dataa(!h2f_WSTRB_6),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_134),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[134] .extended_lut = "off";
defparam \src_data[134] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[134] .shared_arith = "off";

cyclonev_lcell_comb \src_data[138] (
	.dataa(!h2f_WSTRB_10),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_138),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[138] .extended_lut = "off";
defparam \src_data[138] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[138] .shared_arith = "off";

cyclonev_lcell_comb \src_data[142] (
	.dataa(!h2f_WSTRB_14),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_142),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[142] .extended_lut = "off";
defparam \src_data[142] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[142] .shared_arith = "off";

cyclonev_lcell_comb \src_data[146] (
	.dataa(!h2f_ARADDR_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(!out_data_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_146),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[146] .extended_lut = "off";
defparam \src_data[146] .lut_mask = 64'h111F111F111F111F;
defparam \src_data[146] .shared_arith = "off";

cyclonev_lcell_comb \src_data[128] (
	.dataa(!h2f_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_128),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[128] .extended_lut = "off";
defparam \src_data[128] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[128] .shared_arith = "off";

cyclonev_lcell_comb \src_data[132] (
	.dataa(!h2f_WSTRB_4),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_132),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[132] .extended_lut = "off";
defparam \src_data[132] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[132] .shared_arith = "off";

cyclonev_lcell_comb \src_data[136] (
	.dataa(!h2f_WSTRB_8),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_136),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[136] .extended_lut = "off";
defparam \src_data[136] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[136] .shared_arith = "off";

cyclonev_lcell_comb \src_data[140] (
	.dataa(!h2f_WSTRB_12),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_140),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[140] .extended_lut = "off";
defparam \src_data[140] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[140] .shared_arith = "off";

cyclonev_lcell_comb \src_data[129] (
	.dataa(!h2f_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_129),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[129] .extended_lut = "off";
defparam \src_data[129] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[129] .shared_arith = "off";

cyclonev_lcell_comb \src_data[133] (
	.dataa(!h2f_WSTRB_5),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_133),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[133] .extended_lut = "off";
defparam \src_data[133] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[133] .shared_arith = "off";

cyclonev_lcell_comb \src_data[137] (
	.dataa(!h2f_WSTRB_9),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_137),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[137] .extended_lut = "off";
defparam \src_data[137] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[137] .shared_arith = "off";

cyclonev_lcell_comb \src_data[141] (
	.dataa(!h2f_WSTRB_13),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_141),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[141] .extended_lut = "off";
defparam \src_data[141] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[141] .shared_arith = "off";

cyclonev_lcell_comb \src_data[131] (
	.dataa(!h2f_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_131),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[131] .extended_lut = "off";
defparam \src_data[131] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[131] .shared_arith = "off";

cyclonev_lcell_comb \src_data[135] (
	.dataa(!h2f_WSTRB_7),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_135),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[135] .extended_lut = "off";
defparam \src_data[135] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[135] .shared_arith = "off";

cyclonev_lcell_comb \src_data[139] (
	.dataa(!h2f_WSTRB_11),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_139),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[139] .extended_lut = "off";
defparam \src_data[139] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[139] .shared_arith = "off";

cyclonev_lcell_comb \src_data[143] (
	.dataa(!h2f_WSTRB_15),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_143),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[143] .extended_lut = "off";
defparam \src_data[143] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \src_data[143] .shared_arith = "off";

cyclonev_lcell_comb \src_data[184] (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_AWLEN_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(!sop_enable),
	.dataf(!burst_bytecount_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_184),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[184] .extended_lut = "off";
defparam \src_data[184] .lut_mask = 64'h0ACE0A0A0ACE0AFF;
defparam \src_data[184] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!h2f_AWLEN_2),
	.datad(!saved_grant_0),
	.datae(!sop_enable),
	.dataf(!burst_bytecount_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h001E0000001E00FF;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h001E001E001E001E;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!h2f_AWLEN_0),
	.datab(!h2f_AWLEN_1),
	.datac(!saved_grant_0),
	.datad(!sop_enable),
	.datae(!burst_bytecount_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h0600060F0600060F;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h0606060606060606;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[187] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!sop_enable),
	.datad(!burst_bytecount_7),
	.datae(!Add0),
	.dataf(!Add2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_187),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[187] .extended_lut = "off";
defparam \src_data[187] .lut_mask = 64'h0003303355577577;
defparam \src_data[187] .shared_arith = "off";

cyclonev_lcell_comb \src_data[186] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!sop_enable),
	.datad(!burst_bytecount_6),
	.datae(!Add01),
	.dataf(!Add21),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_186),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[186] .extended_lut = "off";
defparam \src_data[186] .lut_mask = 64'h0003303355577577;
defparam \src_data[186] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!h2f_ARLEN_3),
	.datae(!saved_grant_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h0000000100000001;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[188] (
	.dataa(!saved_grant_0),
	.datab(!write_cp_data_188),
	.datac(!src_payload6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_188),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[188] .extended_lut = "off";
defparam \src_data[188] .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \src_data[188] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!h2f_ARLEN_3),
	.datae(!saved_grant_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h000001FE000001FE;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_valid~1 (
	.dataa(!saved_grant_0),
	.datab(!Equal0),
	.datac(!Equal01),
	.datad(!Equal02),
	.datae(!src1_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~1 .extended_lut = "off";
defparam \src_valid~1 .lut_mask = 64'h0000555400005554;
defparam \src_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!saved_grant_0),
	.datad(!LessThan12),
	.datae(!Add42),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h07050F0D07050F0D;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[191]~6 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!saved_grant_1),
	.datad(!\src_data[189]~2_combout ),
	.datae(!Add52),
	.dataf(!\src_data[191]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_191),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[191]~6 .extended_lut = "off";
defparam \src_data[191]~6 .lut_mask = 64'h07050F0D07070F0F;
defparam \src_data[191]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!saved_grant_0),
	.datad(!Selector26),
	.datae(!Add43),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h07050F0D07050F0D;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[192]~7 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!saved_grant_1),
	.datad(!\src_data[189]~2_combout ),
	.datae(!Add53),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_192),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[192]~7 .extended_lut = "off";
defparam \src_data[192]~7 .lut_mask = 64'h07050F0D07050F0D;
defparam \src_data[192]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[193]~8 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!saved_grant_0),
	.datad(!LessThan14),
	.datae(!Add44),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_193),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[193]~8 .extended_lut = "off";
defparam \src_data[193]~8 .lut_mask = 64'h07050F0D07050F0D;
defparam \src_data[193]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[193]~10 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!saved_grant_1),
	.datad(!Add54),
	.datae(!\src_data[193]~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1931),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[193]~10 .extended_lut = "off";
defparam \src_data[193]~10 .lut_mask = 64'h070F050D070F050D;
defparam \src_data[193]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!h2f_ARADDR_4),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h1111111111111111;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[194]~12 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!saved_grant_1),
	.datad(!Add55),
	.datae(!\src_data[194]~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_194),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[194]~12 .extended_lut = "off";
defparam \src_data[194]~12 .lut_mask = 64'h070F050D070F050D;
defparam \src_data[194]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[194]~13 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!saved_grant_0),
	.datad(!LessThan15),
	.datae(!Add45),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1941),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[194]~13 .extended_lut = "off";
defparam \src_data[194]~13 .lut_mask = 64'h07050F0D07050F0D;
defparam \src_data[194]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!h2f_ARADDR_5),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h1111111111111111;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[195]~15 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!saved_grant_1),
	.datad(!Add56),
	.datae(!\src_data[195]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_195),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[195]~15 .extended_lut = "off";
defparam \src_data[195]~15 .lut_mask = 64'h070F050D070F050D;
defparam \src_data[195]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[195]~16 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!saved_grant_0),
	.datad(!LessThan16),
	.datae(!Add46),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1951),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[195]~16 .extended_lut = "off";
defparam \src_data[195]~16 .lut_mask = 64'h07050F0D07050F0D;
defparam \src_data[195]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!h2f_ARADDR_6),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h1111111111111111;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[196]~17 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!saved_grant_0),
	.datad(!Add1),
	.datae(!Add47),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_196),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[196]~17 .extended_lut = "off";
defparam \src_data[196]~17 .lut_mask = 64'h05070D0F05070D0F;
defparam \src_data[196]~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[196]~18 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!saved_grant_1),
	.datad(!Add32),
	.datae(!Add57),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1961),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[196]~18 .extended_lut = "off";
defparam \src_data[196]~18 .lut_mask = 64'h05070D0F05070D0F;
defparam \src_data[196]~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!h2f_ARADDR_7),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h1111111111111111;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[197]~19 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!saved_grant_0),
	.datad(!Add48),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_197),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[197]~19 .extended_lut = "off";
defparam \src_data[197]~19 .lut_mask = 64'h050D050D050D050D;
defparam \src_data[197]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_data[197]~20 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!saved_grant_1),
	.datad(!Add58),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1971),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[197]~20 .extended_lut = "off";
defparam \src_data[197]~20 .lut_mask = 64'h050D050D050D050D;
defparam \src_data[197]~20 .shared_arith = "off";

cyclonev_lcell_comb \src_data[152] (
	.dataa(!h2f_ARADDR_8),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(!out_data_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_152),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[152] .extended_lut = "off";
defparam \src_data[152] .lut_mask = 64'h111F111F111F111F;
defparam \src_data[152] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_0),
	.datab(!out_data_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h1111111111111111;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!h2f_ARADDR_9),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h1111111111111111;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[190]~22 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector7),
	.datad(!\src_data[190]~21_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1901),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[190]~22 .extended_lut = "off";
defparam \src_data[190]~22 .lut_mask = 64'h7530753075307530;
defparam \src_data[190]~22 .shared_arith = "off";

cyclonev_lcell_comb \src_data[189]~24 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector8),
	.datad(!\src_data[189]~23_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1891),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[189]~24 .extended_lut = "off";
defparam \src_data[189]~24 .lut_mask = 64'h7530753075307530;
defparam \src_data[189]~24 .shared_arith = "off";

cyclonev_lcell_comb \src_data[209] (
	.dataa(!h2f_ARID_0),
	.datab(!h2f_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_209),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[209] .extended_lut = "off";
defparam \src_data[209] .lut_mask = 64'h0537053705370537;
defparam \src_data[209] .shared_arith = "off";

cyclonev_lcell_comb \src_data[210] (
	.dataa(!h2f_ARID_1),
	.datab(!h2f_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_210),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[210] .extended_lut = "off";
defparam \src_data[210] .lut_mask = 64'h0537053705370537;
defparam \src_data[210] .shared_arith = "off";

cyclonev_lcell_comb \src_data[211] (
	.dataa(!h2f_ARID_2),
	.datab(!h2f_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_211),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[211] .extended_lut = "off";
defparam \src_data[211] .lut_mask = 64'h0537053705370537;
defparam \src_data[211] .shared_arith = "off";

cyclonev_lcell_comb \src_data[212] (
	.dataa(!h2f_ARID_3),
	.datab(!h2f_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_212),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[212] .extended_lut = "off";
defparam \src_data[212] .lut_mask = 64'h0537053705370537;
defparam \src_data[212] .shared_arith = "off";

cyclonev_lcell_comb \src_data[213] (
	.dataa(!h2f_ARID_4),
	.datab(!h2f_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_213),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[213] .extended_lut = "off";
defparam \src_data[213] .lut_mask = 64'h0537053705370537;
defparam \src_data[213] .shared_arith = "off";

cyclonev_lcell_comb \src_data[214] (
	.dataa(!h2f_ARID_5),
	.datab(!h2f_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_214),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[214] .extended_lut = "off";
defparam \src_data[214] .lut_mask = 64'h0537053705370537;
defparam \src_data[214] .shared_arith = "off";

cyclonev_lcell_comb \src_data[215] (
	.dataa(!h2f_ARID_6),
	.datab(!h2f_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_215),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[215] .extended_lut = "off";
defparam \src_data[215] .lut_mask = 64'h0537053705370537;
defparam \src_data[215] .shared_arith = "off";

cyclonev_lcell_comb \src_data[216] (
	.dataa(!h2f_ARID_7),
	.datab(!h2f_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_216),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[216] .extended_lut = "off";
defparam \src_data[216] .lut_mask = 64'h0537053705370537;
defparam \src_data[216] .shared_arith = "off";

cyclonev_lcell_comb \src_data[217] (
	.dataa(!h2f_ARID_8),
	.datab(!h2f_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_217),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[217] .extended_lut = "off";
defparam \src_data[217] .lut_mask = 64'h0537053705370537;
defparam \src_data[217] .shared_arith = "off";

cyclonev_lcell_comb \src_data[218] (
	.dataa(!h2f_ARID_9),
	.datab(!h2f_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_218),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[218] .extended_lut = "off";
defparam \src_data[218] .lut_mask = 64'h0537053705370537;
defparam \src_data[218] .shared_arith = "off";

cyclonev_lcell_comb \src_data[219] (
	.dataa(!h2f_ARID_10),
	.datab(!h2f_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_219),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[219] .extended_lut = "off";
defparam \src_data[219] .lut_mask = 64'h0537053705370537;
defparam \src_data[219] .shared_arith = "off";

cyclonev_lcell_comb \src_data[220] (
	.dataa(!h2f_ARID_11),
	.datab(!h2f_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_220),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[220] .extended_lut = "off";
defparam \src_data[220] .lut_mask = 64'h0537053705370537;
defparam \src_data[220] .shared_arith = "off";

cyclonev_lcell_comb \src_data[191]~26 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!\src_data[191]~25_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1911),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[191]~26 .extended_lut = "off";
defparam \src_data[191]~26 .lut_mask = 64'h7530753075307530;
defparam \src_data[191]~26 .shared_arith = "off";

cyclonev_lcell_comb \src_data[192]~28 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!\src_data[192]~27_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1921),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[192]~28 .extended_lut = "off";
defparam \src_data[192]~28 .lut_mask = 64'h7530753075307530;
defparam \src_data[192]~28 .shared_arith = "off";

cyclonev_lcell_comb \src_data[193]~31 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!\src_data[193]~29_combout ),
	.datad(!\src_data[193]~30_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1932),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[193]~31 .extended_lut = "off";
defparam \src_data[193]~31 .lut_mask = 64'h7530753075307530;
defparam \src_data[193]~31 .shared_arith = "off";

cyclonev_lcell_comb \src_data[194]~34 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!\src_data[194]~32_combout ),
	.datad(!\src_data[194]~33_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1942),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[194]~34 .extended_lut = "off";
defparam \src_data[194]~34 .lut_mask = 64'h7350735073507350;
defparam \src_data[194]~34 .shared_arith = "off";

cyclonev_lcell_comb \src_data[195]~37 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!\src_data[195]~35_combout ),
	.datad(!\src_data[195]~36_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1952),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[195]~37 .extended_lut = "off";
defparam \src_data[195]~37 .lut_mask = 64'h7350735073507350;
defparam \src_data[195]~37 .shared_arith = "off";

cyclonev_lcell_comb \src_data[196]~40 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!\src_data[196]~38_combout ),
	.datad(!\src_data[196]~39_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1962),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[196]~40 .extended_lut = "off";
defparam \src_data[196]~40 .lut_mask = 64'h7530753075307530;
defparam \src_data[196]~40 .shared_arith = "off";

cyclonev_lcell_comb \src_data[197]~42 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(!\src_data[197]~41_combout ),
	.dataf(!Add58),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1972),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[197]~42 .extended_lut = "off";
defparam \src_data[197]~42 .lut_mask = 64'h05FF05050DFF0D0D;
defparam \src_data[197]~42 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(outclk_wire_0),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!in_ready),
	.datab(!nxt_in_ready),
	.datac(!nxt_in_ready1),
	.datad(!WideOr11),
	.datae(!src_payload_0),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFF00FFA2000000A2;
defparam \update_grant~0 .shared_arith = "off";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!saved_grant_1),
	.datab(!cmd_src_valid_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h1111111111111111;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[190]~0 (
	.dataa(!h2f_ARLEN_3),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(!Add3),
	.datae(!log2ceil),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[190]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[190]~0 .extended_lut = "off";
defparam \src_data[190]~0 .lut_mask = 64'h8000000080000000;
defparam \src_data[190]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[189]~2 (
	.dataa(!h2f_ARLEN_3),
	.datab(!h2f_ARSIZE_2),
	.datac(!Add31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[189]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[189]~2 .extended_lut = "off";
defparam \src_data[189]~2 .lut_mask = 64'h8080808080808080;
defparam \src_data[189]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[189]~3 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!h2f_ARLEN_3),
	.datae(!h2f_ARSIZE_0),
	.dataf(!h2f_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[189]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[189]~3 .extended_lut = "off";
defparam \src_data[189]~3 .lut_mask = 64'h80FF0F0030004000;
defparam \src_data[189]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[191]~5 (
	.dataa(!h2f_ARLEN_0),
	.datab(!h2f_ARLEN_1),
	.datac(!h2f_ARLEN_2),
	.datad(!h2f_ARLEN_3),
	.datae(!h2f_ARSIZE_0),
	.dataf(!h2f_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[191]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[191]~5 .extended_lut = "off";
defparam \src_data[191]~5 .lut_mask = 64'h0F003000400080FF;
defparam \src_data[191]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[193]~9 (
	.dataa(!h2f_ARLEN_3),
	.datab(!h2f_ARSIZE_2),
	.datac(!Add31),
	.datad(!\src_data[189]~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[193]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[193]~9 .extended_lut = "off";
defparam \src_data[193]~9 .lut_mask = 64'h80E880E880E880E8;
defparam \src_data[193]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[194]~11 (
	.dataa(!h2f_ARLEN_3),
	.datab(!h2f_ARSIZE_1),
	.datac(!h2f_ARSIZE_2),
	.datad(!Add3),
	.datae(!log2ceil),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[194]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[194]~11 .extended_lut = "off";
defparam \src_data[194]~11 .lut_mask = 64'hE8A0A080E8A0A080;
defparam \src_data[194]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[195]~14 (
	.dataa(!h2f_ARLEN_3),
	.datab(!h2f_ARSIZE_2),
	.datac(!Add31),
	.datad(!\src_data[191]~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[195]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[195]~14 .extended_lut = "off";
defparam \src_data[195]~14 .lut_mask = 64'hE880E880E880E880;
defparam \src_data[195]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[190]~21 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!Add5),
	.datad(!\src_data[190]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[190]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[190]~21 .extended_lut = "off";
defparam \src_data[190]~21 .lut_mask = 64'h80A280A280A280A2;
defparam \src_data[190]~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[189]~23 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!\src_data[189]~2_combout ),
	.datad(!Add51),
	.datae(!\src_data[189]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[189]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[189]~23 .extended_lut = "off";
defparam \src_data[189]~23 .lut_mask = 64'h88008A0288008A02;
defparam \src_data[189]~23 .shared_arith = "off";

cyclonev_lcell_comb \src_data[191]~25 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!\src_data[189]~2_combout ),
	.datad(!Add52),
	.datae(!\src_data[191]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[191]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[191]~25 .extended_lut = "off";
defparam \src_data[191]~25 .lut_mask = 64'h8A0288008A028800;
defparam \src_data[191]~25 .shared_arith = "off";

cyclonev_lcell_comb \src_data[192]~27 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!\src_data[189]~2_combout ),
	.datad(!Add53),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[192]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[192]~27 .extended_lut = "off";
defparam \src_data[192]~27 .lut_mask = 64'h8A028A028A028A02;
defparam \src_data[192]~27 .shared_arith = "off";

cyclonev_lcell_comb \src_data[193]~29 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!LessThan14),
	.datad(!Add44),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[193]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[193]~29 .extended_lut = "off";
defparam \src_data[193]~29 .lut_mask = 64'h8A028A028A028A02;
defparam \src_data[193]~29 .shared_arith = "off";

cyclonev_lcell_comb \src_data[193]~30 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!Add54),
	.datad(!\src_data[193]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[193]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[193]~30 .extended_lut = "off";
defparam \src_data[193]~30 .lut_mask = 64'h80A280A280A280A2;
defparam \src_data[193]~30 .shared_arith = "off";

cyclonev_lcell_comb \src_data[194]~32 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!Add55),
	.datad(!\src_data[194]~11_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[194]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[194]~32 .extended_lut = "off";
defparam \src_data[194]~32 .lut_mask = 64'h80A280A280A280A2;
defparam \src_data[194]~32 .shared_arith = "off";

cyclonev_lcell_comb \src_data[194]~33 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!LessThan15),
	.datad(!Add45),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[194]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[194]~33 .extended_lut = "off";
defparam \src_data[194]~33 .lut_mask = 64'h8A028A028A028A02;
defparam \src_data[194]~33 .shared_arith = "off";

cyclonev_lcell_comb \src_data[195]~35 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!Add56),
	.datad(!\src_data[195]~14_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[195]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[195]~35 .extended_lut = "off";
defparam \src_data[195]~35 .lut_mask = 64'h80A280A280A280A2;
defparam \src_data[195]~35 .shared_arith = "off";

cyclonev_lcell_comb \src_data[195]~36 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!LessThan16),
	.datad(!Add46),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[195]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[195]~36 .extended_lut = "off";
defparam \src_data[195]~36 .lut_mask = 64'h8A028A028A028A02;
defparam \src_data[195]~36 .shared_arith = "off";

cyclonev_lcell_comb \src_data[196]~38 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!Add1),
	.datad(!Add47),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[196]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[196]~38 .extended_lut = "off";
defparam \src_data[196]~38 .lut_mask = 64'hA820A820A820A820;
defparam \src_data[196]~38 .shared_arith = "off";

cyclonev_lcell_comb \src_data[196]~39 (
	.dataa(!h2f_ARBURST_0),
	.datab(!h2f_ARBURST_1),
	.datac(!Add32),
	.datad(!Add57),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[196]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[196]~39 .extended_lut = "off";
defparam \src_data[196]~39 .lut_mask = 64'hA820A820A820A820;
defparam \src_data[196]~39 .shared_arith = "off";

cyclonev_lcell_comb \src_data[197]~41 (
	.dataa(!h2f_AWBURST_0),
	.datab(!h2f_AWBURST_1),
	.datac(!Add48),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[197]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[197]~41 .extended_lut = "off";
defparam \src_data[197]~41 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \src_data[197]~41 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_arbitrator (
	clk,
	in_ready,
	nxt_in_ready,
	Equal0,
	Equal01,
	Equal02,
	reset,
	Equal03,
	cmd_src_valid_1,
	src1_valid,
	grant_1,
	WideOr1,
	src_payload_0,
	packet_in_progress,
	grant_0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	in_ready;
input 	nxt_in_ready;
input 	Equal0;
input 	Equal01;
input 	Equal02;
input 	reset;
input 	Equal03;
input 	cmd_src_valid_1;
input 	src1_valid;
output 	grant_1;
input 	WideOr1;
input 	src_payload_0;
input 	packet_in_progress;
output 	grant_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!Equal03),
	.datab(!cmd_src_valid_1),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!\top_priority_reg[0]~q ),
	.datae(!src1_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h3303130333031303;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!Equal03),
	.datab(!cmd_src_valid_1),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!\top_priority_reg[0]~q ),
	.datae(!src1_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0000AA080000AA08;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!Equal0),
	.datab(!Equal01),
	.datac(!Equal02),
	.datad(!cmd_src_valid_1),
	.datae(!src1_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFF000100FF000100;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!in_ready),
	.datab(!nxt_in_ready),
	.datac(!WideOr1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hF0F8000800000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module Computer_System_altera_merlin_arbitrator_1 (
	clk,
	Equal0,
	Equal01,
	reset,
	src0_valid,
	update_grant,
	last_cycle,
	grant_0,
	nxt_in_ready,
	nxt_in_ready1,
	src0_valid1,
	sink_ready)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	Equal0;
input 	Equal01;
input 	reset;
input 	src0_valid;
input 	update_grant;
input 	last_cycle;
output 	grant_0;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	src0_valid1;
input 	sink_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!Equal0),
	.datab(!Equal01),
	.datac(!src0_valid),
	.datad(!\top_priority_reg[1]~q ),
	.datae(!\top_priority_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'h0101000101010001;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!nxt_in_ready),
	.datab(!nxt_in_ready1),
	.datac(!sink_ready),
	.datad(!src0_valid1),
	.datae(!update_grant),
	.dataf(!last_cycle),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'h000000FF000700FF;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_router (
	h2f_AWADDR_2,
	h2f_AWADDR_3,
	h2f_AWADDR_4,
	h2f_AWADDR_5,
	h2f_AWADDR_6,
	h2f_AWADDR_7,
	h2f_AWADDR_8,
	h2f_AWADDR_9,
	h2f_AWADDR_10,
	h2f_AWADDR_11,
	h2f_AWADDR_12,
	h2f_AWADDR_13,
	h2f_AWADDR_14,
	h2f_AWADDR_15,
	h2f_AWADDR_16,
	h2f_AWADDR_17,
	h2f_AWADDR_18,
	h2f_AWADDR_19,
	h2f_AWADDR_20,
	h2f_AWADDR_21,
	h2f_AWADDR_22,
	h2f_AWADDR_23,
	h2f_AWADDR_24,
	h2f_AWADDR_25,
	h2f_AWADDR_26,
	h2f_AWADDR_27,
	address_burst_24,
	address_burst_25,
	address_burst_23,
	address_burst_13,
	address_burst_21,
	address_burst_22,
	address_burst_19,
	address_burst_20,
	address_burst_15,
	address_burst_16,
	address_burst_17,
	address_burst_18,
	address_burst_26,
	address_burst_27,
	address_burst_12,
	address_burst_14,
	address_burst_10,
	address_burst_11,
	address_burst_9,
	address_burst_8,
	sop_enable,
	Equal0,
	Equal01,
	address_burst_7,
	address_burst_6,
	address_burst_2,
	address_burst_3,
	address_burst_4,
	address_burst_5,
	Equal02,
	Equal03,
	Equal04)/* synthesis synthesis_greybox=0 */;
input 	h2f_AWADDR_2;
input 	h2f_AWADDR_3;
input 	h2f_AWADDR_4;
input 	h2f_AWADDR_5;
input 	h2f_AWADDR_6;
input 	h2f_AWADDR_7;
input 	h2f_AWADDR_8;
input 	h2f_AWADDR_9;
input 	h2f_AWADDR_10;
input 	h2f_AWADDR_11;
input 	h2f_AWADDR_12;
input 	h2f_AWADDR_13;
input 	h2f_AWADDR_14;
input 	h2f_AWADDR_15;
input 	h2f_AWADDR_16;
input 	h2f_AWADDR_17;
input 	h2f_AWADDR_18;
input 	h2f_AWADDR_19;
input 	h2f_AWADDR_20;
input 	h2f_AWADDR_21;
input 	h2f_AWADDR_22;
input 	h2f_AWADDR_23;
input 	h2f_AWADDR_24;
input 	h2f_AWADDR_25;
input 	h2f_AWADDR_26;
input 	h2f_AWADDR_27;
input 	address_burst_24;
input 	address_burst_25;
input 	address_burst_23;
input 	address_burst_13;
input 	address_burst_21;
input 	address_burst_22;
input 	address_burst_19;
input 	address_burst_20;
input 	address_burst_15;
input 	address_burst_16;
input 	address_burst_17;
input 	address_burst_18;
input 	address_burst_26;
input 	address_burst_27;
input 	address_burst_12;
input 	address_burst_14;
input 	address_burst_10;
input 	address_burst_11;
input 	address_burst_9;
input 	address_burst_8;
input 	sop_enable;
output 	Equal0;
output 	Equal01;
input 	address_burst_7;
input 	address_burst_6;
input 	address_burst_2;
input 	address_burst_3;
input 	address_burst_4;
input 	address_burst_5;
output 	Equal02;
output 	Equal03;
output 	Equal04;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \Equal0~3_combout ;
wire \Equal0~4_combout ;
wire \Equal0~5_combout ;
wire \Equal0~8_combout ;
wire \Equal0~9_combout ;
wire \Equal0~10_combout ;
wire \Equal0~11_combout ;
wire \Equal0~12_combout ;
wire \Equal0~13_combout ;
wire \Equal0~15_combout ;


cyclonev_lcell_comb \Equal0~6 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~1_combout ),
	.datac(!\Equal0~2_combout ),
	.datad(!\Equal0~3_combout ),
	.datae(!\Equal0~4_combout ),
	.dataf(!\Equal0~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~6 .extended_lut = "off";
defparam \Equal0~6 .lut_mask = 64'h0000000000000001;
defparam \Equal0~6 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~7 (
	.dataa(!h2f_AWADDR_26),
	.datab(!h2f_AWADDR_27),
	.datac(!sop_enable),
	.datad(!address_burst_26),
	.datae(!address_burst_27),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal01),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~7 .extended_lut = "off";
defparam \Equal0~7 .lut_mask = 64'h8F8080808F808080;
defparam \Equal0~7 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~14 (
	.dataa(!\Equal0~8_combout ),
	.datab(!\Equal0~9_combout ),
	.datac(!\Equal0~10_combout ),
	.datad(!\Equal0~11_combout ),
	.datae(!\Equal0~12_combout ),
	.dataf(!\Equal0~13_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal02),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~14 .extended_lut = "off";
defparam \Equal0~14 .lut_mask = 64'h0000000000000001;
defparam \Equal0~14 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~16 (
	.dataa(!Equal01),
	.datab(!\Equal0~8_combout ),
	.datac(!\Equal0~9_combout ),
	.datad(!\Equal0~10_combout ),
	.datae(!\Equal0~11_combout ),
	.dataf(!\Equal0~15_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal03),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~16 .extended_lut = "off";
defparam \Equal0~16 .lut_mask = 64'h0000000000000001;
defparam \Equal0~16 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~17 (
	.dataa(!Equal0),
	.datab(!Equal01),
	.datac(!Equal02),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal04),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~17 .extended_lut = "off";
defparam \Equal0~17 .lut_mask = 64'h0101010101010101;
defparam \Equal0~17 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!h2f_AWADDR_24),
	.datab(!h2f_AWADDR_25),
	.datac(!sop_enable),
	.datad(!address_burst_24),
	.datae(!address_burst_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h8F8080808F808080;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!h2f_AWADDR_13),
	.datab(!h2f_AWADDR_23),
	.datac(!sop_enable),
	.datad(!address_burst_23),
	.datae(!address_burst_13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'h8F8080808F808080;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~2 (
	.dataa(!h2f_AWADDR_21),
	.datab(!h2f_AWADDR_22),
	.datac(!sop_enable),
	.datad(!address_burst_21),
	.datae(!address_burst_22),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~2 .extended_lut = "off";
defparam \Equal0~2 .lut_mask = 64'h8F8080808F808080;
defparam \Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~3 (
	.dataa(!h2f_AWADDR_19),
	.datab(!h2f_AWADDR_20),
	.datac(!sop_enable),
	.datad(!address_burst_19),
	.datae(!address_burst_20),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~3 .extended_lut = "off";
defparam \Equal0~3 .lut_mask = 64'h8F8080808F808080;
defparam \Equal0~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~4 (
	.dataa(!h2f_AWADDR_15),
	.datab(!h2f_AWADDR_16),
	.datac(!sop_enable),
	.datad(!address_burst_15),
	.datae(!address_burst_16),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~4 .extended_lut = "off";
defparam \Equal0~4 .lut_mask = 64'h8F8080808F808080;
defparam \Equal0~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~5 (
	.dataa(!h2f_AWADDR_17),
	.datab(!h2f_AWADDR_18),
	.datac(!sop_enable),
	.datad(!address_burst_17),
	.datae(!address_burst_18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~5 .extended_lut = "off";
defparam \Equal0~5 .lut_mask = 64'h8F8080808F808080;
defparam \Equal0~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~8 (
	.dataa(!h2f_AWADDR_12),
	.datab(!h2f_AWADDR_14),
	.datac(!sop_enable),
	.datad(!address_burst_12),
	.datae(!address_burst_14),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~8 .extended_lut = "off";
defparam \Equal0~8 .lut_mask = 64'h8F8080808F808080;
defparam \Equal0~8 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~9 (
	.dataa(!h2f_AWADDR_10),
	.datab(!h2f_AWADDR_11),
	.datac(!sop_enable),
	.datad(!address_burst_10),
	.datae(!address_burst_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~9 .extended_lut = "off";
defparam \Equal0~9 .lut_mask = 64'h8F8080808F808080;
defparam \Equal0~9 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~10 (
	.dataa(!h2f_AWADDR_7),
	.datab(!h2f_AWADDR_9),
	.datac(!sop_enable),
	.datad(!address_burst_7),
	.datae(!address_burst_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~10 .extended_lut = "off";
defparam \Equal0~10 .lut_mask = 64'h8F8080808F808080;
defparam \Equal0~10 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~11 (
	.dataa(!h2f_AWADDR_6),
	.datab(!h2f_AWADDR_8),
	.datac(!sop_enable),
	.datad(!address_burst_6),
	.datae(!address_burst_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~11 .extended_lut = "off";
defparam \Equal0~11 .lut_mask = 64'h8F8080808F808080;
defparam \Equal0~11 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~12 (
	.dataa(!h2f_AWADDR_2),
	.datab(!h2f_AWADDR_3),
	.datac(!sop_enable),
	.datad(!address_burst_2),
	.datae(!address_burst_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~12 .extended_lut = "off";
defparam \Equal0~12 .lut_mask = 64'h8F8080808F808080;
defparam \Equal0~12 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~13 (
	.dataa(!h2f_AWADDR_4),
	.datab(!h2f_AWADDR_5),
	.datac(!sop_enable),
	.datad(!address_burst_4),
	.datae(!address_burst_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~13 .extended_lut = "off";
defparam \Equal0~13 .lut_mask = 64'h8F8080808F808080;
defparam \Equal0~13 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~15 (
	.dataa(!\Equal0~12_combout ),
	.datab(!\Equal0~13_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~15 .extended_lut = "off";
defparam \Equal0~15 .lut_mask = 64'h1111111111111111;
defparam \Equal0~15 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_rsp_demux (
	mem_68_0,
	comb,
	ShiftRight0,
	always10,
	always101,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=0 */;
input 	mem_68_0;
input 	comb;
input 	ShiftRight0;
input 	always10;
input 	always101;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always10),
	.datae(!always101),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'h1111001011110010;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always10),
	.datae(!always101),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h2222002022220020;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_rsp_demux_1 (
	mem_66_0,
	mem_68_0,
	src0_valid)/* synthesis synthesis_greybox=0 */;
input 	mem_66_0;
input 	mem_68_0;
output 	src0_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!mem_66_0),
	.datab(!mem_68_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'h2222222222222222;
defparam \src0_valid~0 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_rsp_mux (
	out_valid,
	src_payload,
	always10,
	src0_valid,
	mem_68_0,
	comb,
	ShiftRight0,
	always101,
	always102,
	src0_valid1,
	WideOr11,
	mem_101_0,
	mem_101_01,
	src_data_209,
	mem_102_0,
	mem_102_01,
	src_data_210,
	mem_103_0,
	mem_103_01,
	src_data_211,
	mem_104_0,
	mem_104_01,
	src_data_212,
	mem_105_0,
	mem_105_01,
	src_data_213,
	mem_106_0,
	mem_106_01,
	src_data_214,
	mem_107_0,
	mem_107_01,
	src_data_215,
	mem_108_0,
	mem_108_01,
	src_data_216,
	mem_109_0,
	mem_109_01,
	src_data_217,
	mem_110_0,
	mem_110_01,
	src_data_218,
	mem_111_0,
	mem_111_01,
	src_data_219,
	mem_112_0,
	mem_112_01,
	src_data_220)/* synthesis synthesis_greybox=0 */;
input 	out_valid;
input 	src_payload;
input 	always10;
input 	src0_valid;
input 	mem_68_0;
input 	comb;
input 	ShiftRight0;
input 	always101;
input 	always102;
input 	src0_valid1;
output 	WideOr11;
input 	mem_101_0;
input 	mem_101_01;
output 	src_data_209;
input 	mem_102_0;
input 	mem_102_01;
output 	src_data_210;
input 	mem_103_0;
input 	mem_103_01;
output 	src_data_211;
input 	mem_104_0;
input 	mem_104_01;
output 	src_data_212;
input 	mem_105_0;
input 	mem_105_01;
output 	src_data_213;
input 	mem_106_0;
input 	mem_106_01;
output 	src_data_214;
input 	mem_107_0;
input 	mem_107_01;
output 	src_data_215;
input 	mem_108_0;
input 	mem_108_01;
output 	src_data_216;
input 	mem_109_0;
input 	mem_109_01;
output 	src_data_217;
input 	mem_110_0;
input 	mem_110_01;
output 	src_data_218;
input 	mem_111_0;
input 	mem_111_01;
output 	src_data_219;
input 	mem_112_0;
input 	mem_112_01;
output 	src_data_220;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_payload~0_combout ;
wire \src_payload~1_combout ;
wire \src_payload~2_combout ;
wire \src_payload~3_combout ;
wire \src_payload~4_combout ;
wire \src_payload~5_combout ;
wire \src_payload~6_combout ;
wire \src_payload~7_combout ;
wire \src_payload~8_combout ;
wire \src_payload~9_combout ;
wire \src_payload~10_combout ;
wire \src_payload~11_combout ;


cyclonev_lcell_comb WideOr1(
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!src0_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h00A2FFFF00A2FFFF;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[209] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~0_combout ),
	.dataf(!mem_101_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_209),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[209] .extended_lut = "off";
defparam \src_data[209] .lut_mask = 64'h0000FFFF00A2FFFF;
defparam \src_data[209] .shared_arith = "off";

cyclonev_lcell_comb \src_data[210] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~1_combout ),
	.dataf(!mem_102_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_210),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[210] .extended_lut = "off";
defparam \src_data[210] .lut_mask = 64'h0000FFFF00A2FFFF;
defparam \src_data[210] .shared_arith = "off";

cyclonev_lcell_comb \src_data[211] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!mem_103_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_211),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[211] .extended_lut = "off";
defparam \src_data[211] .lut_mask = 64'h0000FFFF00A2FFFF;
defparam \src_data[211] .shared_arith = "off";

cyclonev_lcell_comb \src_data[212] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~3_combout ),
	.dataf(!mem_104_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_212),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[212] .extended_lut = "off";
defparam \src_data[212] .lut_mask = 64'h0000FFFF00A2FFFF;
defparam \src_data[212] .shared_arith = "off";

cyclonev_lcell_comb \src_data[213] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~4_combout ),
	.dataf(!mem_105_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_213),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[213] .extended_lut = "off";
defparam \src_data[213] .lut_mask = 64'h0000FFFF00A2FFFF;
defparam \src_data[213] .shared_arith = "off";

cyclonev_lcell_comb \src_data[214] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~5_combout ),
	.dataf(!mem_106_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_214),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[214] .extended_lut = "off";
defparam \src_data[214] .lut_mask = 64'h0000FFFF00A2FFFF;
defparam \src_data[214] .shared_arith = "off";

cyclonev_lcell_comb \src_data[215] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~6_combout ),
	.dataf(!mem_107_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_215),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[215] .extended_lut = "off";
defparam \src_data[215] .lut_mask = 64'h0000FFFF00A2FFFF;
defparam \src_data[215] .shared_arith = "off";

cyclonev_lcell_comb \src_data[216] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~7_combout ),
	.dataf(!mem_108_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_216),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[216] .extended_lut = "off";
defparam \src_data[216] .lut_mask = 64'h0000FFFF00A2FFFF;
defparam \src_data[216] .shared_arith = "off";

cyclonev_lcell_comb \src_data[217] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~8_combout ),
	.dataf(!mem_109_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_217),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[217] .extended_lut = "off";
defparam \src_data[217] .lut_mask = 64'h0000FFFF00A2FFFF;
defparam \src_data[217] .shared_arith = "off";

cyclonev_lcell_comb \src_data[218] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~9_combout ),
	.dataf(!mem_110_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_218),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[218] .extended_lut = "off";
defparam \src_data[218] .lut_mask = 64'h0000FFFF00A2FFFF;
defparam \src_data[218] .shared_arith = "off";

cyclonev_lcell_comb \src_data[219] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~10_combout ),
	.dataf(!mem_111_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_219),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[219] .extended_lut = "off";
defparam \src_data[219] .lut_mask = 64'h0000FFFF00A2FFFF;
defparam \src_data[219] .shared_arith = "off";

cyclonev_lcell_comb \src_data[220] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~11_combout ),
	.dataf(!mem_112_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_220),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[220] .extended_lut = "off";
defparam \src_data[220] .lut_mask = 64'h0000FFFF00A2FFFF;
defparam \src_data[220] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_101_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h0000000011110010;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_102_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h0000000011110010;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_103_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h0000000011110010;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_104_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h0000000011110010;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_105_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h0000000011110010;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_106_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h0000000011110010;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_107_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h0000000011110010;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_108_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h0000000011110010;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_109_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h0000000011110010;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_110_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h0000000011110010;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_111_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h0000000011110010;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!mem_68_0),
	.datab(!comb),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_112_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h0000000011110010;
defparam \src_payload~11 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_0_rsp_mux_1 (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	data_reg_0,
	data_reg_01,
	data_reg_1,
	data_reg_2,
	data_reg_3,
	data_reg_4,
	data_reg_5,
	data_reg_6,
	data_reg_7,
	data_reg_8,
	data_reg_9,
	data_reg_10,
	data_reg_11,
	data_reg_12,
	data_reg_13,
	data_reg_14,
	data_reg_15,
	data_reg_16,
	data_reg_17,
	data_reg_18,
	data_reg_19,
	data_reg_20,
	data_reg_21,
	data_reg_22,
	data_reg_23,
	data_reg_24,
	data_reg_25,
	data_reg_26,
	data_reg_27,
	data_reg_28,
	data_reg_29,
	data_reg_30,
	data_reg_31,
	data_reg_32,
	data_reg_321,
	data_reg_33,
	data_reg_34,
	data_reg_35,
	data_reg_36,
	data_reg_37,
	data_reg_38,
	data_reg_39,
	data_reg_40,
	data_reg_41,
	data_reg_42,
	data_reg_43,
	data_reg_44,
	data_reg_45,
	data_reg_46,
	data_reg_47,
	data_reg_48,
	data_reg_49,
	data_reg_50,
	data_reg_51,
	data_reg_52,
	data_reg_53,
	data_reg_54,
	data_reg_55,
	data_reg_56,
	data_reg_57,
	data_reg_58,
	data_reg_59,
	data_reg_60,
	data_reg_61,
	data_reg_62,
	data_reg_63,
	data_reg_64,
	data_reg_641,
	data_reg_65,
	data_reg_66,
	data_reg_67,
	data_reg_68,
	data_reg_69,
	data_reg_70,
	data_reg_71,
	data_reg_72,
	data_reg_73,
	data_reg_74,
	data_reg_75,
	data_reg_76,
	data_reg_77,
	data_reg_78,
	data_reg_79,
	data_reg_80,
	data_reg_81,
	data_reg_82,
	data_reg_83,
	data_reg_84,
	data_reg_85,
	data_reg_86,
	data_reg_87,
	data_reg_88,
	data_reg_89,
	data_reg_90,
	data_reg_91,
	data_reg_92,
	data_reg_93,
	data_reg_94,
	data_reg_95,
	out_valid,
	comb,
	mem_126_0,
	mem_66_0,
	burst_uncompress_busy,
	last_packet_beat,
	last_packet_beat1,
	last_packet_beat2,
	src_payload,
	mem_38_0,
	source_addr_2,
	mem_39_0,
	source_addr_3,
	always10,
	src0_valid,
	mem_68_0,
	comb1,
	ShiftRight0,
	source_addr_21,
	always101,
	mem_126_01,
	source_addr_31,
	always102,
	src_payload_0,
	src1_valid,
	WideOr11,
	mem_101_0,
	mem_101_01,
	mem_102_0,
	mem_102_01,
	mem_103_0,
	mem_103_01,
	mem_104_0,
	mem_104_01,
	mem_105_0,
	mem_105_01,
	mem_106_0,
	mem_106_01,
	mem_107_0,
	mem_107_01,
	mem_108_0,
	mem_108_01,
	mem_109_0,
	mem_109_01,
	mem_110_0,
	mem_110_01,
	mem_111_0,
	mem_111_01,
	mem_112_0,
	mem_112_01,
	mem_31_0,
	LessThan15,
	ShiftLeft0,
	always4,
	mem_0_0,
	LessThan151,
	src_data_0,
	mem_1_0,
	src_payload1,
	mem_2_0,
	src_data_2,
	mem_3_0,
	src_data_3,
	mem_4_0,
	src_payload2,
	mem_5_0,
	src_data_5,
	mem_6_0,
	src_payload3,
	mem_7_0,
	src_data_7,
	mem_8_0,
	src_payload4,
	mem_9_0,
	src_data_9,
	mem_10_0,
	src_data_10,
	mem_11_0,
	src_data_11,
	mem_12_0,
	src_data_12,
	mem_13_0,
	src_payload5,
	mem_14_0,
	src_data_14,
	mem_15_0,
	src_data_15,
	mem_16_0,
	src_data_16,
	mem_17_0,
	src_payload6,
	mem_18_0,
	src_data_18,
	mem_19_0,
	src_data_19,
	mem_20_0,
	src_payload7,
	mem_21_0,
	src_data_21,
	mem_22_0,
	src_payload8,
	mem_23_0,
	src_data_23,
	mem_24_0,
	src_payload9,
	mem_25_0,
	src_data_25,
	mem_26_0,
	src_data_26,
	mem_27_0,
	src_data_27,
	mem_28_0,
	src_data_28,
	mem_29_0,
	src_payload10,
	mem_30_0,
	src_data_30,
	mem_31_01,
	src_data_31,
	ShiftLeft01,
	src_data_32,
	src_payload11,
	src_data_34,
	src_data_35,
	src_payload12,
	src_data_37,
	src_payload13,
	src_data_39,
	src_payload14,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_payload15,
	src_data_46,
	src_data_47,
	src_data_48,
	src_payload16,
	src_data_50,
	src_data_51,
	src_payload17,
	src_data_53,
	src_payload18,
	src_data_55,
	src_payload19,
	src_data_57,
	src_data_58,
	src_data_59,
	src_data_60,
	src_payload20,
	src_data_62,
	src_data_63,
	ShiftLeft02,
	src_data_64,
	src_payload21,
	src_data_66,
	src_data_67,
	src_payload22,
	src_data_69,
	src_payload23,
	src_data_71,
	src_payload24,
	src_data_73,
	src_data_74,
	src_data_75,
	src_data_76,
	src_payload25,
	src_data_78,
	src_data_79,
	src_data_80,
	src_payload26,
	src_data_82,
	src_data_83,
	src_payload27,
	src_data_85,
	src_payload28,
	src_data_87,
	src_payload29,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_payload30,
	src_data_94,
	src_data_95,
	src_data_96,
	out_data_1,
	src_payload31,
	src_data_98,
	src_data_99,
	out_data_4,
	src_payload32,
	src_data_101,
	out_data_6,
	src_payload33,
	src_data_103,
	out_data_8,
	src_payload34,
	src_data_105,
	src_data_106,
	src_data_107,
	src_data_108,
	out_data_13,
	src_payload35,
	src_data_110,
	src_data_111,
	src_data_112,
	out_data_17,
	src_payload36,
	src_data_114,
	src_data_115,
	out_data_20,
	src_payload37,
	src_data_117,
	out_data_22,
	src_payload38,
	src_data_119,
	out_data_24,
	src_payload39,
	src_data_121,
	src_data_122,
	src_data_123,
	src_data_124,
	out_data_29,
	src_payload40,
	src_data_126,
	src_data_127,
	src_data_209,
	src_data_210,
	src_data_211,
	src_data_212,
	src_data_213,
	src_data_214,
	src_data_215,
	src_data_216,
	src_data_217,
	src_data_218,
	src_data_219,
	src_data_220,
	src_payload41)/* synthesis synthesis_greybox=0 */;
input 	q_b_0;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	q_b_8;
input 	q_b_9;
input 	q_b_10;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_20;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_24;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_28;
input 	q_b_29;
input 	q_b_30;
input 	q_b_31;
input 	data_reg_0;
input 	data_reg_01;
input 	data_reg_1;
input 	data_reg_2;
input 	data_reg_3;
input 	data_reg_4;
input 	data_reg_5;
input 	data_reg_6;
input 	data_reg_7;
input 	data_reg_8;
input 	data_reg_9;
input 	data_reg_10;
input 	data_reg_11;
input 	data_reg_12;
input 	data_reg_13;
input 	data_reg_14;
input 	data_reg_15;
input 	data_reg_16;
input 	data_reg_17;
input 	data_reg_18;
input 	data_reg_19;
input 	data_reg_20;
input 	data_reg_21;
input 	data_reg_22;
input 	data_reg_23;
input 	data_reg_24;
input 	data_reg_25;
input 	data_reg_26;
input 	data_reg_27;
input 	data_reg_28;
input 	data_reg_29;
input 	data_reg_30;
input 	data_reg_31;
input 	data_reg_32;
input 	data_reg_321;
input 	data_reg_33;
input 	data_reg_34;
input 	data_reg_35;
input 	data_reg_36;
input 	data_reg_37;
input 	data_reg_38;
input 	data_reg_39;
input 	data_reg_40;
input 	data_reg_41;
input 	data_reg_42;
input 	data_reg_43;
input 	data_reg_44;
input 	data_reg_45;
input 	data_reg_46;
input 	data_reg_47;
input 	data_reg_48;
input 	data_reg_49;
input 	data_reg_50;
input 	data_reg_51;
input 	data_reg_52;
input 	data_reg_53;
input 	data_reg_54;
input 	data_reg_55;
input 	data_reg_56;
input 	data_reg_57;
input 	data_reg_58;
input 	data_reg_59;
input 	data_reg_60;
input 	data_reg_61;
input 	data_reg_62;
input 	data_reg_63;
input 	data_reg_64;
input 	data_reg_641;
input 	data_reg_65;
input 	data_reg_66;
input 	data_reg_67;
input 	data_reg_68;
input 	data_reg_69;
input 	data_reg_70;
input 	data_reg_71;
input 	data_reg_72;
input 	data_reg_73;
input 	data_reg_74;
input 	data_reg_75;
input 	data_reg_76;
input 	data_reg_77;
input 	data_reg_78;
input 	data_reg_79;
input 	data_reg_80;
input 	data_reg_81;
input 	data_reg_82;
input 	data_reg_83;
input 	data_reg_84;
input 	data_reg_85;
input 	data_reg_86;
input 	data_reg_87;
input 	data_reg_88;
input 	data_reg_89;
input 	data_reg_90;
input 	data_reg_91;
input 	data_reg_92;
input 	data_reg_93;
input 	data_reg_94;
input 	data_reg_95;
input 	out_valid;
input 	comb;
input 	mem_126_0;
input 	mem_66_0;
input 	burst_uncompress_busy;
input 	last_packet_beat;
input 	last_packet_beat1;
input 	last_packet_beat2;
output 	src_payload;
input 	mem_38_0;
input 	source_addr_2;
input 	mem_39_0;
input 	source_addr_3;
input 	always10;
input 	src0_valid;
input 	mem_68_0;
input 	comb1;
input 	ShiftRight0;
input 	source_addr_21;
input 	always101;
input 	mem_126_01;
input 	source_addr_31;
input 	always102;
output 	src_payload_0;
input 	src1_valid;
output 	WideOr11;
input 	mem_101_0;
input 	mem_101_01;
input 	mem_102_0;
input 	mem_102_01;
input 	mem_103_0;
input 	mem_103_01;
input 	mem_104_0;
input 	mem_104_01;
input 	mem_105_0;
input 	mem_105_01;
input 	mem_106_0;
input 	mem_106_01;
input 	mem_107_0;
input 	mem_107_01;
input 	mem_108_0;
input 	mem_108_01;
input 	mem_109_0;
input 	mem_109_01;
input 	mem_110_0;
input 	mem_110_01;
input 	mem_111_0;
input 	mem_111_01;
input 	mem_112_0;
input 	mem_112_01;
input 	mem_31_0;
input 	LessThan15;
input 	ShiftLeft0;
input 	always4;
input 	mem_0_0;
input 	LessThan151;
output 	src_data_0;
input 	mem_1_0;
output 	src_payload1;
input 	mem_2_0;
output 	src_data_2;
input 	mem_3_0;
output 	src_data_3;
input 	mem_4_0;
output 	src_payload2;
input 	mem_5_0;
output 	src_data_5;
input 	mem_6_0;
output 	src_payload3;
input 	mem_7_0;
output 	src_data_7;
input 	mem_8_0;
output 	src_payload4;
input 	mem_9_0;
output 	src_data_9;
input 	mem_10_0;
output 	src_data_10;
input 	mem_11_0;
output 	src_data_11;
input 	mem_12_0;
output 	src_data_12;
input 	mem_13_0;
output 	src_payload5;
input 	mem_14_0;
output 	src_data_14;
input 	mem_15_0;
output 	src_data_15;
input 	mem_16_0;
output 	src_data_16;
input 	mem_17_0;
output 	src_payload6;
input 	mem_18_0;
output 	src_data_18;
input 	mem_19_0;
output 	src_data_19;
input 	mem_20_0;
output 	src_payload7;
input 	mem_21_0;
output 	src_data_21;
input 	mem_22_0;
output 	src_payload8;
input 	mem_23_0;
output 	src_data_23;
input 	mem_24_0;
output 	src_payload9;
input 	mem_25_0;
output 	src_data_25;
input 	mem_26_0;
output 	src_data_26;
input 	mem_27_0;
output 	src_data_27;
input 	mem_28_0;
output 	src_data_28;
input 	mem_29_0;
output 	src_payload10;
input 	mem_30_0;
output 	src_data_30;
input 	mem_31_01;
output 	src_data_31;
input 	ShiftLeft01;
output 	src_data_32;
output 	src_payload11;
output 	src_data_34;
output 	src_data_35;
output 	src_payload12;
output 	src_data_37;
output 	src_payload13;
output 	src_data_39;
output 	src_payload14;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_payload15;
output 	src_data_46;
output 	src_data_47;
output 	src_data_48;
output 	src_payload16;
output 	src_data_50;
output 	src_data_51;
output 	src_payload17;
output 	src_data_53;
output 	src_payload18;
output 	src_data_55;
output 	src_payload19;
output 	src_data_57;
output 	src_data_58;
output 	src_data_59;
output 	src_data_60;
output 	src_payload20;
output 	src_data_62;
output 	src_data_63;
input 	ShiftLeft02;
output 	src_data_64;
output 	src_payload21;
output 	src_data_66;
output 	src_data_67;
output 	src_payload22;
output 	src_data_69;
output 	src_payload23;
output 	src_data_71;
output 	src_payload24;
output 	src_data_73;
output 	src_data_74;
output 	src_data_75;
output 	src_data_76;
output 	src_payload25;
output 	src_data_78;
output 	src_data_79;
output 	src_data_80;
output 	src_payload26;
output 	src_data_82;
output 	src_data_83;
output 	src_payload27;
output 	src_data_85;
output 	src_payload28;
output 	src_data_87;
output 	src_payload29;
output 	src_data_89;
output 	src_data_90;
output 	src_data_91;
output 	src_data_92;
output 	src_payload30;
output 	src_data_94;
output 	src_data_95;
output 	src_data_96;
input 	out_data_1;
output 	src_payload31;
output 	src_data_98;
output 	src_data_99;
input 	out_data_4;
output 	src_payload32;
output 	src_data_101;
input 	out_data_6;
output 	src_payload33;
output 	src_data_103;
input 	out_data_8;
output 	src_payload34;
output 	src_data_105;
output 	src_data_106;
output 	src_data_107;
output 	src_data_108;
input 	out_data_13;
output 	src_payload35;
output 	src_data_110;
output 	src_data_111;
output 	src_data_112;
input 	out_data_17;
output 	src_payload36;
output 	src_data_114;
output 	src_data_115;
input 	out_data_20;
output 	src_payload37;
output 	src_data_117;
input 	out_data_22;
output 	src_payload38;
output 	src_data_119;
input 	out_data_24;
output 	src_payload39;
output 	src_data_121;
output 	src_data_122;
output 	src_data_123;
output 	src_data_124;
input 	out_data_29;
output 	src_payload40;
output 	src_data_126;
output 	src_data_127;
output 	src_data_209;
output 	src_data_210;
output 	src_data_211;
output 	src_data_212;
output 	src_data_213;
output 	src_data_214;
output 	src_data_215;
output 	src_data_216;
output 	src_data_217;
output 	src_data_218;
output 	src_data_219;
output 	src_data_220;
output 	src_payload41;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_payload~1_combout ;
wire \src_payload~2_combout ;
wire \src_data[0]~0_combout ;
wire \src_payload~3_combout ;
wire \src_data[2]~2_combout ;
wire \src_data[3]~4_combout ;
wire \src_payload~5_combout ;
wire \src_data[5]~6_combout ;
wire \src_payload~7_combout ;
wire \src_data[7]~8_combout ;
wire \src_payload~9_combout ;
wire \src_data[9]~10_combout ;
wire \src_data[10]~12_combout ;
wire \src_data[11]~14_combout ;
wire \src_data[12]~16_combout ;
wire \src_payload~11_combout ;
wire \src_data[14]~18_combout ;
wire \src_data[15]~20_combout ;
wire \src_data[16]~22_combout ;
wire \src_payload~13_combout ;
wire \src_data[18]~24_combout ;
wire \src_data[19]~26_combout ;
wire \src_payload~15_combout ;
wire \src_data[21]~28_combout ;
wire \src_payload~17_combout ;
wire \src_data[23]~30_combout ;
wire \src_payload~19_combout ;
wire \src_data[25]~32_combout ;
wire \src_data[26]~34_combout ;
wire \src_data[27]~36_combout ;
wire \src_data[28]~38_combout ;
wire \src_payload~21_combout ;
wire \src_data[30]~40_combout ;
wire \src_data[31]~42_combout ;
wire \src_payload~23_combout ;
wire \src_payload~24_combout ;
wire \src_data[32]~44_combout ;
wire \src_payload~25_combout ;
wire \src_data[34]~46_combout ;
wire \src_data[35]~48_combout ;
wire \src_payload~27_combout ;
wire \src_data[37]~50_combout ;
wire \src_payload~29_combout ;
wire \src_data[39]~52_combout ;
wire \src_payload~31_combout ;
wire \src_data[41]~54_combout ;
wire \src_data[42]~56_combout ;
wire \src_data[43]~58_combout ;
wire \src_data[44]~60_combout ;
wire \src_payload~33_combout ;
wire \src_data[46]~62_combout ;
wire \src_data[47]~64_combout ;
wire \src_data[48]~66_combout ;
wire \src_payload~35_combout ;
wire \src_data[50]~68_combout ;
wire \src_data[51]~70_combout ;
wire \src_payload~37_combout ;
wire \src_data[53]~72_combout ;
wire \src_payload~39_combout ;
wire \src_data[55]~74_combout ;
wire \src_payload~41_combout ;
wire \src_data[57]~76_combout ;
wire \src_data[58]~78_combout ;
wire \src_data[59]~80_combout ;
wire \src_data[60]~82_combout ;
wire \src_payload~43_combout ;
wire \src_data[62]~84_combout ;
wire \src_data[63]~86_combout ;
wire \src_payload~45_combout ;
wire \src_payload~46_combout ;
wire \src_data[64]~88_combout ;
wire \src_payload~47_combout ;
wire \src_data[66]~90_combout ;
wire \src_data[67]~92_combout ;
wire \src_payload~49_combout ;
wire \src_data[69]~94_combout ;
wire \src_payload~51_combout ;
wire \src_data[71]~96_combout ;
wire \src_payload~53_combout ;
wire \src_data[73]~98_combout ;
wire \src_data[74]~100_combout ;
wire \src_data[75]~102_combout ;
wire \src_data[76]~104_combout ;
wire \src_payload~55_combout ;
wire \src_data[78]~106_combout ;
wire \src_data[79]~108_combout ;
wire \src_data[80]~110_combout ;
wire \src_payload~57_combout ;
wire \src_data[82]~112_combout ;
wire \src_data[83]~114_combout ;
wire \src_payload~59_combout ;
wire \src_data[85]~116_combout ;
wire \src_payload~61_combout ;
wire \src_data[87]~118_combout ;
wire \src_payload~63_combout ;
wire \src_data[89]~120_combout ;
wire \src_data[90]~122_combout ;
wire \src_data[91]~124_combout ;
wire \src_data[92]~126_combout ;
wire \src_payload~65_combout ;
wire \src_data[94]~128_combout ;
wire \src_data[95]~130_combout ;
wire \src_payload~67_combout ;
wire \src_payload~68_combout ;
wire \src_payload~69_combout ;
wire \src_payload~70_combout ;
wire \src_payload~81_combout ;
wire \src_payload~82_combout ;
wire \src_payload~83_combout ;
wire \src_payload~84_combout ;
wire \src_payload~85_combout ;
wire \src_payload~86_combout ;
wire \src_payload~87_combout ;
wire \src_payload~88_combout ;
wire \src_payload~89_combout ;
wire \src_payload~90_combout ;
wire \src_payload~91_combout ;
wire \src_payload~92_combout ;


cyclonev_lcell_comb \src_payload~0 (
	.dataa(!comb),
	.datab(!mem_126_0),
	.datac(!mem_66_0),
	.datad(!last_packet_beat),
	.datae(!last_packet_beat1),
	.dataf(!last_packet_beat2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h3030303131313131;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(gnd),
	.datad(!src0_valid),
	.datae(!src_payload41),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h2200FFFF2200FFFF;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!src1_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hA200FFFFA200FFFF;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~1 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~1 .extended_lut = "off";
defparam \src_data[0]~1 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~3 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[2]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~3 .extended_lut = "off";
defparam \src_data[2]~3 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[2]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~5 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[3]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~5 .extended_lut = "off";
defparam \src_data[3]~5 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~7 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[5]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~7 .extended_lut = "off";
defparam \src_data[5]~7 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[5]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~9 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[7]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~9 .extended_lut = "off";
defparam \src_data[7]~9 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[7]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~11 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[9]~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~11 .extended_lut = "off";
defparam \src_data[9]~11 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[9]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[10]~13 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[10]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10]~13 .extended_lut = "off";
defparam \src_data[10]~13 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[10]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[11]~15 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[11]~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11]~15 .extended_lut = "off";
defparam \src_data[11]~15 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[11]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[12]~17 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[12]~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12]~17 .extended_lut = "off";
defparam \src_data[12]~17 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[12]~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[14]~19 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[14]~18_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14]~19 .extended_lut = "off";
defparam \src_data[14]~19 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[14]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_data[15]~21 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[15]~20_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15]~21 .extended_lut = "off";
defparam \src_data[15]~21 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[15]~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[16]~23 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[16]~22_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16]~23 .extended_lut = "off";
defparam \src_data[16]~23 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[16]~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~13_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[18]~25 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[18]~24_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18]~25 .extended_lut = "off";
defparam \src_data[18]~25 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[18]~25 .shared_arith = "off";

cyclonev_lcell_comb \src_data[19]~27 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[19]~26_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19]~27 .extended_lut = "off";
defparam \src_data[19]~27 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[19]~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[21]~29 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[21]~28_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21]~29 .extended_lut = "off";
defparam \src_data[21]~29 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[21]~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~17_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_data[23]~31 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[23]~30_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23]~31 .extended_lut = "off";
defparam \src_data[23]~31 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[23]~31 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_data[25]~33 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[25]~32_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25]~33 .extended_lut = "off";
defparam \src_data[25]~33 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[25]~33 .shared_arith = "off";

cyclonev_lcell_comb \src_data[26]~35 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[26]~34_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26]~35 .extended_lut = "off";
defparam \src_data[26]~35 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[26]~35 .shared_arith = "off";

cyclonev_lcell_comb \src_data[27]~37 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[27]~36_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27]~37 .extended_lut = "off";
defparam \src_data[27]~37 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[27]~37 .shared_arith = "off";

cyclonev_lcell_comb \src_data[28]~39 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[28]~38_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28]~39 .extended_lut = "off";
defparam \src_data[28]~39 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[28]~39 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_data[30]~41 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[30]~40_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30]~41 .extended_lut = "off";
defparam \src_data[30]~41 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[30]~41 .shared_arith = "off";

cyclonev_lcell_comb \src_data[31]~43 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~2_combout ),
	.dataf(!\src_data[31]~42_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31]~43 .extended_lut = "off";
defparam \src_data[31]~43 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[31]~43 .shared_arith = "off";

cyclonev_lcell_comb \src_data[32]~45 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[32]~44_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32]~45 .extended_lut = "off";
defparam \src_data[32]~45 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[32]~45 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34]~47 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[34]~46_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34]~47 .extended_lut = "off";
defparam \src_data[34]~47 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[34]~47 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35]~49 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[35]~48_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35]~49 .extended_lut = "off";
defparam \src_data[35]~49 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[35]~49 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~27_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_data[37]~51 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[37]~50_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_37),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[37]~51 .extended_lut = "off";
defparam \src_data[37]~51 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[37]~51 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~29_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_data[39]~53 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[39]~52_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39]~53 .extended_lut = "off";
defparam \src_data[39]~53 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[39]~53 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~31_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \src_data[41]~55 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[41]~54_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41]~55 .extended_lut = "off";
defparam \src_data[41]~55 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[41]~55 .shared_arith = "off";

cyclonev_lcell_comb \src_data[42]~57 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[42]~56_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42]~57 .extended_lut = "off";
defparam \src_data[42]~57 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[42]~57 .shared_arith = "off";

cyclonev_lcell_comb \src_data[43]~59 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[43]~58_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43]~59 .extended_lut = "off";
defparam \src_data[43]~59 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[43]~59 .shared_arith = "off";

cyclonev_lcell_comb \src_data[44]~61 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[44]~60_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44]~61 .extended_lut = "off";
defparam \src_data[44]~61 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[44]~61 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~34 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~33_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~34 .extended_lut = "off";
defparam \src_payload~34 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~34 .shared_arith = "off";

cyclonev_lcell_comb \src_data[46]~63 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[46]~62_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46]~63 .extended_lut = "off";
defparam \src_data[46]~63 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[46]~63 .shared_arith = "off";

cyclonev_lcell_comb \src_data[47]~65 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[47]~64_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_47),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[47]~65 .extended_lut = "off";
defparam \src_data[47]~65 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[47]~65 .shared_arith = "off";

cyclonev_lcell_comb \src_data[48]~67 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[48]~66_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_48),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[48]~67 .extended_lut = "off";
defparam \src_data[48]~67 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[48]~67 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~36 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~35_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~36 .extended_lut = "off";
defparam \src_payload~36 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~36 .shared_arith = "off";

cyclonev_lcell_comb \src_data[50]~69 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[50]~68_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_50),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[50]~69 .extended_lut = "off";
defparam \src_data[50]~69 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[50]~69 .shared_arith = "off";

cyclonev_lcell_comb \src_data[51]~71 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[51]~70_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_51),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[51]~71 .extended_lut = "off";
defparam \src_data[51]~71 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[51]~71 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~38 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~37_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~38 .extended_lut = "off";
defparam \src_payload~38 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~38 .shared_arith = "off";

cyclonev_lcell_comb \src_data[53]~73 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[53]~72_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_53),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[53]~73 .extended_lut = "off";
defparam \src_data[53]~73 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[53]~73 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~40 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~39_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~40 .extended_lut = "off";
defparam \src_payload~40 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~40 .shared_arith = "off";

cyclonev_lcell_comb \src_data[55]~75 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[55]~74_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_55),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[55]~75 .extended_lut = "off";
defparam \src_data[55]~75 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[55]~75 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~42 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~41_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~42 .extended_lut = "off";
defparam \src_payload~42 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~42 .shared_arith = "off";

cyclonev_lcell_comb \src_data[57]~77 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[57]~76_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_57),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[57]~77 .extended_lut = "off";
defparam \src_data[57]~77 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[57]~77 .shared_arith = "off";

cyclonev_lcell_comb \src_data[58]~79 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[58]~78_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_58),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[58]~79 .extended_lut = "off";
defparam \src_data[58]~79 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[58]~79 .shared_arith = "off";

cyclonev_lcell_comb \src_data[59]~81 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[59]~80_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_59),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[59]~81 .extended_lut = "off";
defparam \src_data[59]~81 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[59]~81 .shared_arith = "off";

cyclonev_lcell_comb \src_data[60]~83 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[60]~82_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_60),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[60]~83 .extended_lut = "off";
defparam \src_data[60]~83 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[60]~83 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~44 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~43_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~44 .extended_lut = "off";
defparam \src_payload~44 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~44 .shared_arith = "off";

cyclonev_lcell_comb \src_data[62]~85 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[62]~84_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_62),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[62]~85 .extended_lut = "off";
defparam \src_data[62]~85 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[62]~85 .shared_arith = "off";

cyclonev_lcell_comb \src_data[63]~87 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~24_combout ),
	.dataf(!\src_data[63]~86_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_63),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[63]~87 .extended_lut = "off";
defparam \src_data[63]~87 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[63]~87 .shared_arith = "off";

cyclonev_lcell_comb \src_data[64]~89 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[64]~88_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_64),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[64]~89 .extended_lut = "off";
defparam \src_data[64]~89 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[64]~89 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~48 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~47_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~48 .extended_lut = "off";
defparam \src_payload~48 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~48 .shared_arith = "off";

cyclonev_lcell_comb \src_data[66]~91 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[66]~90_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_66),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[66]~91 .extended_lut = "off";
defparam \src_data[66]~91 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[66]~91 .shared_arith = "off";

cyclonev_lcell_comb \src_data[67]~93 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[67]~92_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_67),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[67]~93 .extended_lut = "off";
defparam \src_data[67]~93 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[67]~93 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~50 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~49_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~50 .extended_lut = "off";
defparam \src_payload~50 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~50 .shared_arith = "off";

cyclonev_lcell_comb \src_data[69]~95 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[69]~94_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_69),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[69]~95 .extended_lut = "off";
defparam \src_data[69]~95 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[69]~95 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~52 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~51_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~52 .extended_lut = "off";
defparam \src_payload~52 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~52 .shared_arith = "off";

cyclonev_lcell_comb \src_data[71]~97 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[71]~96_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_71),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71]~97 .extended_lut = "off";
defparam \src_data[71]~97 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[71]~97 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~54 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~53_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~54 .extended_lut = "off";
defparam \src_payload~54 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~54 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~99 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[73]~98_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_73),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~99 .extended_lut = "off";
defparam \src_data[73]~99 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[73]~99 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~101 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[74]~100_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_74),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~101 .extended_lut = "off";
defparam \src_data[74]~101 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[74]~101 .shared_arith = "off";

cyclonev_lcell_comb \src_data[75]~103 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[75]~102_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_75),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[75]~103 .extended_lut = "off";
defparam \src_data[75]~103 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[75]~103 .shared_arith = "off";

cyclonev_lcell_comb \src_data[76]~105 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[76]~104_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_76),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[76]~105 .extended_lut = "off";
defparam \src_data[76]~105 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[76]~105 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~56 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~55_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~56 .extended_lut = "off";
defparam \src_payload~56 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~56 .shared_arith = "off";

cyclonev_lcell_comb \src_data[78]~107 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[78]~106_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_78),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[78]~107 .extended_lut = "off";
defparam \src_data[78]~107 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[78]~107 .shared_arith = "off";

cyclonev_lcell_comb \src_data[79]~109 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[79]~108_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79]~109 .extended_lut = "off";
defparam \src_data[79]~109 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[79]~109 .shared_arith = "off";

cyclonev_lcell_comb \src_data[80]~111 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[80]~110_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_80),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[80]~111 .extended_lut = "off";
defparam \src_data[80]~111 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[80]~111 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~58 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~57_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~58 .extended_lut = "off";
defparam \src_payload~58 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~58 .shared_arith = "off";

cyclonev_lcell_comb \src_data[82]~113 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[82]~112_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_82),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[82]~113 .extended_lut = "off";
defparam \src_data[82]~113 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[82]~113 .shared_arith = "off";

cyclonev_lcell_comb \src_data[83]~115 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[83]~114_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_83),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[83]~115 .extended_lut = "off";
defparam \src_data[83]~115 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[83]~115 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~60 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~59_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~60 .extended_lut = "off";
defparam \src_payload~60 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~60 .shared_arith = "off";

cyclonev_lcell_comb \src_data[85]~117 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[85]~116_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_85),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[85]~117 .extended_lut = "off";
defparam \src_data[85]~117 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[85]~117 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~62 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~61_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~62 .extended_lut = "off";
defparam \src_payload~62 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~62 .shared_arith = "off";

cyclonev_lcell_comb \src_data[87]~119 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[87]~118_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_87),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[87]~119 .extended_lut = "off";
defparam \src_data[87]~119 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[87]~119 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~64 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~63_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~64 .extended_lut = "off";
defparam \src_payload~64 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~64 .shared_arith = "off";

cyclonev_lcell_comb \src_data[89]~121 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[89]~120_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_89),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[89]~121 .extended_lut = "off";
defparam \src_data[89]~121 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[89]~121 .shared_arith = "off";

cyclonev_lcell_comb \src_data[90]~123 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[90]~122_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_90),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[90]~123 .extended_lut = "off";
defparam \src_data[90]~123 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[90]~123 .shared_arith = "off";

cyclonev_lcell_comb \src_data[91]~125 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[91]~124_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_91),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[91]~125 .extended_lut = "off";
defparam \src_data[91]~125 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[91]~125 .shared_arith = "off";

cyclonev_lcell_comb \src_data[92]~127 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[92]~126_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_92),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92]~127 .extended_lut = "off";
defparam \src_data[92]~127 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[92]~127 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~66 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~65_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~66 .extended_lut = "off";
defparam \src_payload~66 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~66 .shared_arith = "off";

cyclonev_lcell_comb \src_data[94]~129 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[94]~128_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_94),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94]~129 .extended_lut = "off";
defparam \src_data[94]~129 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[94]~129 .shared_arith = "off";

cyclonev_lcell_comb \src_data[95]~131 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~46_combout ),
	.dataf(!\src_data[95]~130_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_95),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95]~131 .extended_lut = "off";
defparam \src_data[95]~131 .lut_mask = 64'h0000FFFFA200FFFF;
defparam \src_data[95]~131 .shared_arith = "off";

cyclonev_lcell_comb \src_data[96] (
	.dataa(!q_b_0),
	.datab(!always4),
	.datac(!mem_0_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_96),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96] .extended_lut = "off";
defparam \src_data[96] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[96] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~71 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!out_data_1),
	.dataf(!\src_payload~67_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~71 .extended_lut = "off";
defparam \src_payload~71 .lut_mask = 64'h000000000000A200;
defparam \src_payload~71 .shared_arith = "off";

cyclonev_lcell_comb \src_data[98] (
	.dataa(!q_b_2),
	.datab(!always4),
	.datac(!mem_2_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_98),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98] .extended_lut = "off";
defparam \src_data[98] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[98] .shared_arith = "off";

cyclonev_lcell_comb \src_data[99] (
	.dataa(!q_b_3),
	.datab(!always4),
	.datac(!mem_3_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_99),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99] .extended_lut = "off";
defparam \src_data[99] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[99] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~72 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!out_data_4),
	.dataf(!\src_payload~67_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~72 .extended_lut = "off";
defparam \src_payload~72 .lut_mask = 64'h000000000000A200;
defparam \src_payload~72 .shared_arith = "off";

cyclonev_lcell_comb \src_data[101] (
	.dataa(!q_b_5),
	.datab(!always4),
	.datac(!mem_5_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_101),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[101] .extended_lut = "off";
defparam \src_data[101] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[101] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~73 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!out_data_6),
	.dataf(!\src_payload~67_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~73 .extended_lut = "off";
defparam \src_payload~73 .lut_mask = 64'h000000000000A200;
defparam \src_payload~73 .shared_arith = "off";

cyclonev_lcell_comb \src_data[103] (
	.dataa(!q_b_7),
	.datab(!always4),
	.datac(!mem_7_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_103),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[103] .extended_lut = "off";
defparam \src_data[103] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[103] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~74 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!out_data_8),
	.dataf(!\src_payload~67_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~74 .extended_lut = "off";
defparam \src_payload~74 .lut_mask = 64'h000000000000A200;
defparam \src_payload~74 .shared_arith = "off";

cyclonev_lcell_comb \src_data[105] (
	.dataa(!q_b_9),
	.datab(!always4),
	.datac(!mem_9_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_105),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[105] .extended_lut = "off";
defparam \src_data[105] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[105] .shared_arith = "off";

cyclonev_lcell_comb \src_data[106] (
	.dataa(!q_b_10),
	.datab(!always4),
	.datac(!mem_10_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_106),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[106] .extended_lut = "off";
defparam \src_data[106] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[106] .shared_arith = "off";

cyclonev_lcell_comb \src_data[107] (
	.dataa(!q_b_11),
	.datab(!always4),
	.datac(!mem_11_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_107),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[107] .extended_lut = "off";
defparam \src_data[107] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[107] .shared_arith = "off";

cyclonev_lcell_comb \src_data[108] (
	.dataa(!q_b_12),
	.datab(!always4),
	.datac(!mem_12_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_108),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[108] .extended_lut = "off";
defparam \src_data[108] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[108] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~75 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!out_data_13),
	.dataf(!\src_payload~67_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~75 .extended_lut = "off";
defparam \src_payload~75 .lut_mask = 64'h000000000000A200;
defparam \src_payload~75 .shared_arith = "off";

cyclonev_lcell_comb \src_data[110] (
	.dataa(!q_b_14),
	.datab(!always4),
	.datac(!mem_14_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_110),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[110] .extended_lut = "off";
defparam \src_data[110] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[110] .shared_arith = "off";

cyclonev_lcell_comb \src_data[111] (
	.dataa(!q_b_15),
	.datab(!always4),
	.datac(!mem_15_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_111),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[111] .extended_lut = "off";
defparam \src_data[111] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[111] .shared_arith = "off";

cyclonev_lcell_comb \src_data[112] (
	.dataa(!q_b_16),
	.datab(!always4),
	.datac(!mem_16_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_112),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[112] .extended_lut = "off";
defparam \src_data[112] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[112] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~76 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!out_data_17),
	.dataf(!\src_payload~67_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload36),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~76 .extended_lut = "off";
defparam \src_payload~76 .lut_mask = 64'h000000000000A200;
defparam \src_payload~76 .shared_arith = "off";

cyclonev_lcell_comb \src_data[114] (
	.dataa(!q_b_18),
	.datab(!always4),
	.datac(!mem_18_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_114),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[114] .extended_lut = "off";
defparam \src_data[114] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[114] .shared_arith = "off";

cyclonev_lcell_comb \src_data[115] (
	.dataa(!q_b_19),
	.datab(!always4),
	.datac(!mem_19_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_115),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[115] .extended_lut = "off";
defparam \src_data[115] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[115] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~77 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!out_data_20),
	.dataf(!\src_payload~67_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload37),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~77 .extended_lut = "off";
defparam \src_payload~77 .lut_mask = 64'h000000000000A200;
defparam \src_payload~77 .shared_arith = "off";

cyclonev_lcell_comb \src_data[117] (
	.dataa(!q_b_21),
	.datab(!always4),
	.datac(!mem_21_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_117),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[117] .extended_lut = "off";
defparam \src_data[117] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[117] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~78 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!out_data_22),
	.dataf(!\src_payload~67_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~78 .extended_lut = "off";
defparam \src_payload~78 .lut_mask = 64'h000000000000A200;
defparam \src_payload~78 .shared_arith = "off";

cyclonev_lcell_comb \src_data[119] (
	.dataa(!q_b_23),
	.datab(!always4),
	.datac(!mem_23_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_119),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[119] .extended_lut = "off";
defparam \src_data[119] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[119] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~79 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!out_data_24),
	.dataf(!\src_payload~67_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~79 .extended_lut = "off";
defparam \src_payload~79 .lut_mask = 64'h000000000000A200;
defparam \src_payload~79 .shared_arith = "off";

cyclonev_lcell_comb \src_data[121] (
	.dataa(!q_b_25),
	.datab(!always4),
	.datac(!mem_25_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_121),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[121] .extended_lut = "off";
defparam \src_data[121] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[121] .shared_arith = "off";

cyclonev_lcell_comb \src_data[122] (
	.dataa(!q_b_26),
	.datab(!always4),
	.datac(!mem_26_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_122),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[122] .extended_lut = "off";
defparam \src_data[122] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[122] .shared_arith = "off";

cyclonev_lcell_comb \src_data[123] (
	.dataa(!q_b_27),
	.datab(!always4),
	.datac(!mem_27_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_123),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[123] .extended_lut = "off";
defparam \src_data[123] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[123] .shared_arith = "off";

cyclonev_lcell_comb \src_data[124] (
	.dataa(!q_b_28),
	.datab(!always4),
	.datac(!mem_28_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_124),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[124] .extended_lut = "off";
defparam \src_data[124] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[124] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~80 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!out_data_29),
	.dataf(!\src_payload~67_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~80 .extended_lut = "off";
defparam \src_payload~80 .lut_mask = 64'h000000000000A200;
defparam \src_payload~80 .shared_arith = "off";

cyclonev_lcell_comb \src_data[126] (
	.dataa(!q_b_30),
	.datab(!always4),
	.datac(!mem_30_0),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_126),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[126] .extended_lut = "off";
defparam \src_data[126] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[126] .shared_arith = "off";

cyclonev_lcell_comb \src_data[127] (
	.dataa(!q_b_31),
	.datab(!always4),
	.datac(!mem_31_01),
	.datad(!\src_payload~68_combout ),
	.datae(!\src_payload~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_127),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[127] .extended_lut = "off";
defparam \src_data[127] .lut_mask = 64'h001DFFFF001DFFFF;
defparam \src_data[127] .shared_arith = "off";

cyclonev_lcell_comb \src_data[209] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!mem_101_01),
	.dataf(!\src_payload~81_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_209),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[209] .extended_lut = "off";
defparam \src_data[209] .lut_mask = 64'h0000A200FFFFFFFF;
defparam \src_data[209] .shared_arith = "off";

cyclonev_lcell_comb \src_data[210] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!mem_102_01),
	.dataf(!\src_payload~82_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_210),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[210] .extended_lut = "off";
defparam \src_data[210] .lut_mask = 64'h0000A200FFFFFFFF;
defparam \src_data[210] .shared_arith = "off";

cyclonev_lcell_comb \src_data[211] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!mem_103_01),
	.dataf(!\src_payload~83_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_211),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[211] .extended_lut = "off";
defparam \src_data[211] .lut_mask = 64'h0000A200FFFFFFFF;
defparam \src_data[211] .shared_arith = "off";

cyclonev_lcell_comb \src_data[212] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!mem_104_01),
	.dataf(!\src_payload~84_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_212),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[212] .extended_lut = "off";
defparam \src_data[212] .lut_mask = 64'h0000A200FFFFFFFF;
defparam \src_data[212] .shared_arith = "off";

cyclonev_lcell_comb \src_data[213] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!mem_105_01),
	.dataf(!\src_payload~85_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_213),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[213] .extended_lut = "off";
defparam \src_data[213] .lut_mask = 64'h0000A200FFFFFFFF;
defparam \src_data[213] .shared_arith = "off";

cyclonev_lcell_comb \src_data[214] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!mem_106_01),
	.dataf(!\src_payload~86_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_214),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[214] .extended_lut = "off";
defparam \src_data[214] .lut_mask = 64'h0000A200FFFFFFFF;
defparam \src_data[214] .shared_arith = "off";

cyclonev_lcell_comb \src_data[215] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!mem_107_01),
	.dataf(!\src_payload~87_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_215),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[215] .extended_lut = "off";
defparam \src_data[215] .lut_mask = 64'h0000A200FFFFFFFF;
defparam \src_data[215] .shared_arith = "off";

cyclonev_lcell_comb \src_data[216] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!mem_108_01),
	.dataf(!\src_payload~88_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_216),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[216] .extended_lut = "off";
defparam \src_data[216] .lut_mask = 64'h0000A200FFFFFFFF;
defparam \src_data[216] .shared_arith = "off";

cyclonev_lcell_comb \src_data[217] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!mem_109_01),
	.dataf(!\src_payload~89_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_217),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[217] .extended_lut = "off";
defparam \src_data[217] .lut_mask = 64'h0000A200FFFFFFFF;
defparam \src_data[217] .shared_arith = "off";

cyclonev_lcell_comb \src_data[218] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!mem_110_01),
	.dataf(!\src_payload~90_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_218),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[218] .extended_lut = "off";
defparam \src_data[218] .lut_mask = 64'h0000A200FFFFFFFF;
defparam \src_data[218] .shared_arith = "off";

cyclonev_lcell_comb \src_data[219] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!mem_111_01),
	.dataf(!\src_payload~91_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_219),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[219] .extended_lut = "off";
defparam \src_data[219] .lut_mask = 64'h0000A200FFFFFFFF;
defparam \src_data[219] .shared_arith = "off";

cyclonev_lcell_comb \src_data[220] (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!mem_112_01),
	.dataf(!\src_payload~92_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_220),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[220] .extended_lut = "off";
defparam \src_data[220] .lut_mask = 64'h0000A200FFFFFFFF;
defparam \src_data[220] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~93 (
	.dataa(!comb1),
	.datab(!mem_126_01),
	.datac(!mem_68_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~93 .extended_lut = "off";
defparam \src_payload~93 .lut_mask = 64'h1010101010101010;
defparam \src_payload~93 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!source_addr_21),
	.datab(!source_addr_31),
	.datac(!mem_31_0),
	.datad(!data_reg_0),
	.datae(!LessThan15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h01FF010101FF0101;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!\src_payload~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h0000000022220020;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~0 (
	.dataa(!q_b_0),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!mem_0_0),
	.datae(!data_reg_01),
	.dataf(!LessThan151),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~0 .extended_lut = "off";
defparam \src_data[0]~0 .lut_mask = 64'h0131FFFF01310131;
defparam \src_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!q_b_1),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_1_0),
	.dataf(!data_reg_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h01013131FF01FF31;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~2 (
	.dataa(!q_b_2),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_2_0),
	.dataf(!data_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~2 .extended_lut = "off";
defparam \src_data[2]~2 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~4 (
	.dataa(!q_b_3),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_3_0),
	.dataf(!data_reg_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~4 .extended_lut = "off";
defparam \src_data[3]~4 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!q_b_4),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_4_0),
	.dataf(!data_reg_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h01013131FF01FF31;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~6 (
	.dataa(!q_b_5),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_5_0),
	.dataf(!data_reg_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~6 .extended_lut = "off";
defparam \src_data[5]~6 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[5]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!q_b_6),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_6_0),
	.dataf(!data_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h01013131FF01FF31;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~8 (
	.dataa(!q_b_7),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_7_0),
	.dataf(!data_reg_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~8 .extended_lut = "off";
defparam \src_data[7]~8 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[7]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!q_b_8),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_8_0),
	.dataf(!data_reg_8),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h01013131FF01FF31;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~10 (
	.dataa(!q_b_9),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_9_0),
	.dataf(!data_reg_9),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[9]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~10 .extended_lut = "off";
defparam \src_data[9]~10 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[9]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[10]~12 (
	.dataa(!q_b_10),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_10_0),
	.dataf(!data_reg_10),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[10]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10]~12 .extended_lut = "off";
defparam \src_data[10]~12 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[10]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[11]~14 (
	.dataa(!q_b_11),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_11_0),
	.dataf(!data_reg_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[11]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11]~14 .extended_lut = "off";
defparam \src_data[11]~14 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[11]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[12]~16 (
	.dataa(!q_b_12),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_12_0),
	.dataf(!data_reg_12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[12]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12]~16 .extended_lut = "off";
defparam \src_data[12]~16 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[12]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!q_b_13),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_13_0),
	.dataf(!data_reg_13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h01013131FF01FF31;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[14]~18 (
	.dataa(!q_b_14),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_14_0),
	.dataf(!data_reg_14),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[14]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14]~18 .extended_lut = "off";
defparam \src_data[14]~18 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[14]~18 .shared_arith = "off";

cyclonev_lcell_comb \src_data[15]~20 (
	.dataa(!q_b_15),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_15_0),
	.dataf(!data_reg_15),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[15]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15]~20 .extended_lut = "off";
defparam \src_data[15]~20 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[15]~20 .shared_arith = "off";

cyclonev_lcell_comb \src_data[16]~22 (
	.dataa(!q_b_16),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_16_0),
	.dataf(!data_reg_16),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[16]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16]~22 .extended_lut = "off";
defparam \src_data[16]~22 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[16]~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!q_b_17),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_17_0),
	.dataf(!data_reg_17),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h01013131FF01FF31;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[18]~24 (
	.dataa(!q_b_18),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_18_0),
	.dataf(!data_reg_18),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[18]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18]~24 .extended_lut = "off";
defparam \src_data[18]~24 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[18]~24 .shared_arith = "off";

cyclonev_lcell_comb \src_data[19]~26 (
	.dataa(!q_b_19),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_19_0),
	.dataf(!data_reg_19),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[19]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19]~26 .extended_lut = "off";
defparam \src_data[19]~26 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[19]~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!q_b_20),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_20_0),
	.dataf(!data_reg_20),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h01013131FF01FF31;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[21]~28 (
	.dataa(!q_b_21),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_21_0),
	.dataf(!data_reg_21),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[21]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21]~28 .extended_lut = "off";
defparam \src_data[21]~28 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[21]~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!q_b_22),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_22_0),
	.dataf(!data_reg_22),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h01013131FF01FF31;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[23]~30 (
	.dataa(!q_b_23),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_23_0),
	.dataf(!data_reg_23),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[23]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23]~30 .extended_lut = "off";
defparam \src_data[23]~30 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[23]~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!q_b_24),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_24_0),
	.dataf(!data_reg_24),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h01013131FF01FF31;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_data[25]~32 (
	.dataa(!q_b_25),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_25_0),
	.dataf(!data_reg_25),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[25]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25]~32 .extended_lut = "off";
defparam \src_data[25]~32 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[25]~32 .shared_arith = "off";

cyclonev_lcell_comb \src_data[26]~34 (
	.dataa(!q_b_26),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_26_0),
	.dataf(!data_reg_26),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[26]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26]~34 .extended_lut = "off";
defparam \src_data[26]~34 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[26]~34 .shared_arith = "off";

cyclonev_lcell_comb \src_data[27]~36 (
	.dataa(!q_b_27),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_27_0),
	.dataf(!data_reg_27),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[27]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27]~36 .extended_lut = "off";
defparam \src_data[27]~36 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[27]~36 .shared_arith = "off";

cyclonev_lcell_comb \src_data[28]~38 (
	.dataa(!q_b_28),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_28_0),
	.dataf(!data_reg_28),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[28]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28]~38 .extended_lut = "off";
defparam \src_data[28]~38 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[28]~38 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!q_b_29),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_29_0),
	.dataf(!data_reg_29),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h01013131FF01FF31;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[30]~40 (
	.dataa(!q_b_30),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_30_0),
	.dataf(!data_reg_30),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[30]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30]~40 .extended_lut = "off";
defparam \src_data[30]~40 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[30]~40 .shared_arith = "off";

cyclonev_lcell_comb \src_data[31]~42 (
	.dataa(!q_b_31),
	.datab(!ShiftLeft0),
	.datac(!always4),
	.datad(!LessThan151),
	.datae(!mem_31_01),
	.dataf(!data_reg_31),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[31]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31]~42 .extended_lut = "off";
defparam \src_data[31]~42 .lut_mask = 64'h01013131FF01FF31;
defparam \src_data[31]~42 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!source_addr_21),
	.datab(!source_addr_31),
	.datac(!mem_31_0),
	.datad(!LessThan15),
	.datae(!data_reg_32),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h0202FF020202FF02;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!\src_payload~23_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h0000000022220020;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_data[32]~44 (
	.dataa(!q_b_0),
	.datab(!always4),
	.datac(!mem_0_0),
	.datad(!LessThan151),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_321),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[32]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32]~44 .extended_lut = "off";
defparam \src_data[32]~44 .lut_mask = 64'h00001D1DFF00FF1D;
defparam \src_data[32]~44 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!q_b_1),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_1_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_33),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34]~46 (
	.dataa(!q_b_2),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_2_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_34),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[34]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34]~46 .extended_lut = "off";
defparam \src_data[34]~46 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[34]~46 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35]~48 (
	.dataa(!q_b_3),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_3_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_35),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[35]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35]~48 .extended_lut = "off";
defparam \src_data[35]~48 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[35]~48 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!q_b_4),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_4_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_36),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_data[37]~50 (
	.dataa(!q_b_5),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_5_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_37),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[37]~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[37]~50 .extended_lut = "off";
defparam \src_data[37]~50 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[37]~50 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!q_b_6),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_6_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_38),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_data[39]~52 (
	.dataa(!q_b_7),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_7_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_39),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[39]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39]~52 .extended_lut = "off";
defparam \src_data[39]~52 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[39]~52 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!q_b_8),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_8_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_40),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_data[41]~54 (
	.dataa(!q_b_9),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_9_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_41),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[41]~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41]~54 .extended_lut = "off";
defparam \src_data[41]~54 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[41]~54 .shared_arith = "off";

cyclonev_lcell_comb \src_data[42]~56 (
	.dataa(!q_b_10),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_10_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_42),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[42]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42]~56 .extended_lut = "off";
defparam \src_data[42]~56 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[42]~56 .shared_arith = "off";

cyclonev_lcell_comb \src_data[43]~58 (
	.dataa(!q_b_11),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_11_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_43),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[43]~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43]~58 .extended_lut = "off";
defparam \src_data[43]~58 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[43]~58 .shared_arith = "off";

cyclonev_lcell_comb \src_data[44]~60 (
	.dataa(!q_b_12),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_12_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_44),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[44]~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44]~60 .extended_lut = "off";
defparam \src_data[44]~60 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[44]~60 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~33 (
	.dataa(!q_b_13),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_13_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_45),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~33 .extended_lut = "off";
defparam \src_payload~33 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~33 .shared_arith = "off";

cyclonev_lcell_comb \src_data[46]~62 (
	.dataa(!q_b_14),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_14_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_46),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[46]~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46]~62 .extended_lut = "off";
defparam \src_data[46]~62 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[46]~62 .shared_arith = "off";

cyclonev_lcell_comb \src_data[47]~64 (
	.dataa(!q_b_15),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_15_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_47),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[47]~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[47]~64 .extended_lut = "off";
defparam \src_data[47]~64 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[47]~64 .shared_arith = "off";

cyclonev_lcell_comb \src_data[48]~66 (
	.dataa(!q_b_16),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_16_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_48),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[48]~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[48]~66 .extended_lut = "off";
defparam \src_data[48]~66 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[48]~66 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~35 (
	.dataa(!q_b_17),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_17_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_49),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~35 .extended_lut = "off";
defparam \src_payload~35 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~35 .shared_arith = "off";

cyclonev_lcell_comb \src_data[50]~68 (
	.dataa(!q_b_18),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_18_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_50),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[50]~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[50]~68 .extended_lut = "off";
defparam \src_data[50]~68 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[50]~68 .shared_arith = "off";

cyclonev_lcell_comb \src_data[51]~70 (
	.dataa(!q_b_19),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_19_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_51),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[51]~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[51]~70 .extended_lut = "off";
defparam \src_data[51]~70 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[51]~70 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~37 (
	.dataa(!q_b_20),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_20_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_52),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~37 .extended_lut = "off";
defparam \src_payload~37 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~37 .shared_arith = "off";

cyclonev_lcell_comb \src_data[53]~72 (
	.dataa(!q_b_21),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_21_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_53),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[53]~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[53]~72 .extended_lut = "off";
defparam \src_data[53]~72 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[53]~72 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~39 (
	.dataa(!q_b_22),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_22_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_54),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~39 .extended_lut = "off";
defparam \src_payload~39 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~39 .shared_arith = "off";

cyclonev_lcell_comb \src_data[55]~74 (
	.dataa(!q_b_23),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_23_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_55),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[55]~74_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[55]~74 .extended_lut = "off";
defparam \src_data[55]~74 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[55]~74 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~41 (
	.dataa(!q_b_24),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_24_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_56),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~41 .extended_lut = "off";
defparam \src_payload~41 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~41 .shared_arith = "off";

cyclonev_lcell_comb \src_data[57]~76 (
	.dataa(!q_b_25),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_25_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_57),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[57]~76_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[57]~76 .extended_lut = "off";
defparam \src_data[57]~76 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[57]~76 .shared_arith = "off";

cyclonev_lcell_comb \src_data[58]~78 (
	.dataa(!q_b_26),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_26_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_58),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[58]~78_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[58]~78 .extended_lut = "off";
defparam \src_data[58]~78 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[58]~78 .shared_arith = "off";

cyclonev_lcell_comb \src_data[59]~80 (
	.dataa(!q_b_27),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_27_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_59),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[59]~80_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[59]~80 .extended_lut = "off";
defparam \src_data[59]~80 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[59]~80 .shared_arith = "off";

cyclonev_lcell_comb \src_data[60]~82 (
	.dataa(!q_b_28),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_28_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_60),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[60]~82_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[60]~82 .extended_lut = "off";
defparam \src_data[60]~82 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[60]~82 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~43 (
	.dataa(!q_b_29),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_29_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_61),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~43 .extended_lut = "off";
defparam \src_payload~43 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~43 .shared_arith = "off";

cyclonev_lcell_comb \src_data[62]~84 (
	.dataa(!q_b_30),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_30_0),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_62),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[62]~84_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[62]~84 .extended_lut = "off";
defparam \src_data[62]~84 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[62]~84 .shared_arith = "off";

cyclonev_lcell_comb \src_data[63]~86 (
	.dataa(!q_b_31),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_31_01),
	.datae(!ShiftLeft01),
	.dataf(!data_reg_63),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[63]~86_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[63]~86 .extended_lut = "off";
defparam \src_data[63]~86 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[63]~86 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~45 (
	.dataa(!source_addr_21),
	.datab(!source_addr_31),
	.datac(!mem_31_0),
	.datad(!LessThan15),
	.datae(!data_reg_64),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~45 .extended_lut = "off";
defparam \src_payload~45 .lut_mask = 64'h0404FF040404FF04;
defparam \src_payload~45 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~46 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!\src_payload~45_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~46 .extended_lut = "off";
defparam \src_payload~46 .lut_mask = 64'h0000000022220020;
defparam \src_payload~46 .shared_arith = "off";

cyclonev_lcell_comb \src_data[64]~88 (
	.dataa(!q_b_0),
	.datab(!always4),
	.datac(!mem_0_0),
	.datad(!LessThan151),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_641),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[64]~88_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[64]~88 .extended_lut = "off";
defparam \src_data[64]~88 .lut_mask = 64'h00001D1DFF00FF1D;
defparam \src_data[64]~88 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~47 (
	.dataa(!q_b_1),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_1_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_65),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~47 .extended_lut = "off";
defparam \src_payload~47 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~47 .shared_arith = "off";

cyclonev_lcell_comb \src_data[66]~90 (
	.dataa(!q_b_2),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_2_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_66),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[66]~90_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[66]~90 .extended_lut = "off";
defparam \src_data[66]~90 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[66]~90 .shared_arith = "off";

cyclonev_lcell_comb \src_data[67]~92 (
	.dataa(!q_b_3),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_3_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_67),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[67]~92_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[67]~92 .extended_lut = "off";
defparam \src_data[67]~92 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[67]~92 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~49 (
	.dataa(!q_b_4),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_4_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_68),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~49 .extended_lut = "off";
defparam \src_payload~49 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~49 .shared_arith = "off";

cyclonev_lcell_comb \src_data[69]~94 (
	.dataa(!q_b_5),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_5_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_69),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[69]~94_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[69]~94 .extended_lut = "off";
defparam \src_data[69]~94 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[69]~94 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~51 (
	.dataa(!q_b_6),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_6_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_70),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~51 .extended_lut = "off";
defparam \src_payload~51 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~51 .shared_arith = "off";

cyclonev_lcell_comb \src_data[71]~96 (
	.dataa(!q_b_7),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_7_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_71),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[71]~96_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71]~96 .extended_lut = "off";
defparam \src_data[71]~96 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[71]~96 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~53 (
	.dataa(!q_b_8),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_8_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_72),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~53 .extended_lut = "off";
defparam \src_payload~53 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~53 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~98 (
	.dataa(!q_b_9),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_9_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_73),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[73]~98_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~98 .extended_lut = "off";
defparam \src_data[73]~98 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[73]~98 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~100 (
	.dataa(!q_b_10),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_10_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_74),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[74]~100_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~100 .extended_lut = "off";
defparam \src_data[74]~100 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[74]~100 .shared_arith = "off";

cyclonev_lcell_comb \src_data[75]~102 (
	.dataa(!q_b_11),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_11_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_75),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[75]~102_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[75]~102 .extended_lut = "off";
defparam \src_data[75]~102 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[75]~102 .shared_arith = "off";

cyclonev_lcell_comb \src_data[76]~104 (
	.dataa(!q_b_12),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_12_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_76),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[76]~104_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[76]~104 .extended_lut = "off";
defparam \src_data[76]~104 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[76]~104 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~55 (
	.dataa(!q_b_13),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_13_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_77),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~55 .extended_lut = "off";
defparam \src_payload~55 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~55 .shared_arith = "off";

cyclonev_lcell_comb \src_data[78]~106 (
	.dataa(!q_b_14),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_14_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_78),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[78]~106_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[78]~106 .extended_lut = "off";
defparam \src_data[78]~106 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[78]~106 .shared_arith = "off";

cyclonev_lcell_comb \src_data[79]~108 (
	.dataa(!q_b_15),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_15_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_79),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[79]~108_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79]~108 .extended_lut = "off";
defparam \src_data[79]~108 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[79]~108 .shared_arith = "off";

cyclonev_lcell_comb \src_data[80]~110 (
	.dataa(!q_b_16),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_16_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_80),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[80]~110_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[80]~110 .extended_lut = "off";
defparam \src_data[80]~110 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[80]~110 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~57 (
	.dataa(!q_b_17),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_17_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_81),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~57 .extended_lut = "off";
defparam \src_payload~57 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~57 .shared_arith = "off";

cyclonev_lcell_comb \src_data[82]~112 (
	.dataa(!q_b_18),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_18_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_82),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[82]~112_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[82]~112 .extended_lut = "off";
defparam \src_data[82]~112 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[82]~112 .shared_arith = "off";

cyclonev_lcell_comb \src_data[83]~114 (
	.dataa(!q_b_19),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_19_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_83),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[83]~114_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[83]~114 .extended_lut = "off";
defparam \src_data[83]~114 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[83]~114 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~59 (
	.dataa(!q_b_20),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_20_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_84),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~59 .extended_lut = "off";
defparam \src_payload~59 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~59 .shared_arith = "off";

cyclonev_lcell_comb \src_data[85]~116 (
	.dataa(!q_b_21),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_21_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_85),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[85]~116_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[85]~116 .extended_lut = "off";
defparam \src_data[85]~116 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[85]~116 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~61 (
	.dataa(!q_b_22),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_22_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_86),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~61 .extended_lut = "off";
defparam \src_payload~61 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~61 .shared_arith = "off";

cyclonev_lcell_comb \src_data[87]~118 (
	.dataa(!q_b_23),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_23_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_87),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[87]~118_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[87]~118 .extended_lut = "off";
defparam \src_data[87]~118 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[87]~118 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~63 (
	.dataa(!q_b_24),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_24_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_88),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~63 .extended_lut = "off";
defparam \src_payload~63 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~63 .shared_arith = "off";

cyclonev_lcell_comb \src_data[89]~120 (
	.dataa(!q_b_25),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_25_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_89),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[89]~120_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[89]~120 .extended_lut = "off";
defparam \src_data[89]~120 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[89]~120 .shared_arith = "off";

cyclonev_lcell_comb \src_data[90]~122 (
	.dataa(!q_b_26),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_26_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_90),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[90]~122_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[90]~122 .extended_lut = "off";
defparam \src_data[90]~122 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[90]~122 .shared_arith = "off";

cyclonev_lcell_comb \src_data[91]~124 (
	.dataa(!q_b_27),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_27_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_91),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[91]~124_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[91]~124 .extended_lut = "off";
defparam \src_data[91]~124 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[91]~124 .shared_arith = "off";

cyclonev_lcell_comb \src_data[92]~126 (
	.dataa(!q_b_28),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_28_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_92),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[92]~126_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92]~126 .extended_lut = "off";
defparam \src_data[92]~126 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[92]~126 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~65 (
	.dataa(!q_b_29),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_29_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_93),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~65 .extended_lut = "off";
defparam \src_payload~65 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_payload~65 .shared_arith = "off";

cyclonev_lcell_comb \src_data[94]~128 (
	.dataa(!q_b_30),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_30_0),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_94),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[94]~128_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94]~128 .extended_lut = "off";
defparam \src_data[94]~128 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[94]~128 .shared_arith = "off";

cyclonev_lcell_comb \src_data[95]~130 (
	.dataa(!q_b_31),
	.datab(!always4),
	.datac(!LessThan151),
	.datad(!mem_31_01),
	.datae(!ShiftLeft02),
	.dataf(!data_reg_95),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[95]~130_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95]~130 .extended_lut = "off";
defparam \src_data[95]~130 .lut_mask = 64'h000011DDF0F0F1FD;
defparam \src_data[95]~130 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~67 (
	.dataa(!comb),
	.datab(!burst_uncompress_busy),
	.datac(!mem_38_0),
	.datad(!source_addr_2),
	.datae(!mem_39_0),
	.dataf(!source_addr_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~67 .extended_lut = "off";
defparam \src_payload~67 .lut_mask = 64'hBB00BF0400000404;
defparam \src_payload~67 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~68 (
	.dataa(!out_valid),
	.datab(!src_payload),
	.datac(!always10),
	.datad(!src0_valid),
	.datae(!\src_payload~67_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~68 .extended_lut = "off";
defparam \src_payload~68 .lut_mask = 64'h0000A2000000A200;
defparam \src_payload~68 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~69 (
	.dataa(!source_addr_21),
	.datab(!source_addr_31),
	.datac(!mem_31_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~69 .extended_lut = "off";
defparam \src_payload~69 .lut_mask = 64'h0808080808080808;
defparam \src_payload~69 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~70 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!\src_payload~69_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~70 .extended_lut = "off";
defparam \src_payload~70 .lut_mask = 64'h0000000022220020;
defparam \src_payload~70 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~81 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_101_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~81_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~81 .extended_lut = "off";
defparam \src_payload~81 .lut_mask = 64'h0000000022220020;
defparam \src_payload~81 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~82 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_102_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~82_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~82 .extended_lut = "off";
defparam \src_payload~82 .lut_mask = 64'h0000000022220020;
defparam \src_payload~82 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~83 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_103_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~83_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~83 .extended_lut = "off";
defparam \src_payload~83 .lut_mask = 64'h0000000022220020;
defparam \src_payload~83 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~84 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_104_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~84_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~84 .extended_lut = "off";
defparam \src_payload~84 .lut_mask = 64'h0000000022220020;
defparam \src_payload~84 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~85 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_105_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~85_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~85 .extended_lut = "off";
defparam \src_payload~85 .lut_mask = 64'h0000000022220020;
defparam \src_payload~85 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~86 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_106_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~86_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~86 .extended_lut = "off";
defparam \src_payload~86 .lut_mask = 64'h0000000022220020;
defparam \src_payload~86 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~87 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_107_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~87_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~87 .extended_lut = "off";
defparam \src_payload~87 .lut_mask = 64'h0000000022220020;
defparam \src_payload~87 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~88 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_108_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~88_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~88 .extended_lut = "off";
defparam \src_payload~88 .lut_mask = 64'h0000000022220020;
defparam \src_payload~88 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~89 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_109_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~89_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~89 .extended_lut = "off";
defparam \src_payload~89 .lut_mask = 64'h0000000022220020;
defparam \src_payload~89 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~90 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_110_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~90_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~90 .extended_lut = "off";
defparam \src_payload~90 .lut_mask = 64'h0000000022220020;
defparam \src_payload~90 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~91 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_111_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~91_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~91 .extended_lut = "off";
defparam \src_payload~91 .lut_mask = 64'h0000000022220020;
defparam \src_payload~91 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~92 (
	.dataa(!mem_68_0),
	.datab(!comb1),
	.datac(!ShiftRight0),
	.datad(!always101),
	.datae(!always102),
	.dataf(!mem_112_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~92_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~92 .extended_lut = "off";
defparam \src_payload~92 .lut_mask = 64'h0000000022220020;
defparam \src_payload~92 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_1 (
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	outclk_wire_0,
	in_ready_hold,
	wait_latency_counter_0,
	wait_latency_counter_1,
	sink1_ready,
	ARM_A9_HPS_h2f_lw_axi_master_awready,
	src0_valid,
	source_endofpacket,
	src1_valid,
	ARM_A9_HPS_h2f_lw_axi_master_wready,
	mem_88_0,
	mem_89_0,
	mem_90_0,
	mem_91_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	r_sync_rst,
	m0_write,
	m0_read,
	wrclk_control_slave_readdata_0,
	wrclk_control_slave_readdata_1,
	wrclk_control_slave_readdata_2,
	wrclk_control_slave_readdata_3,
	wrclk_control_slave_readdata_4,
	wrclk_control_slave_readdata_5,
	wrclk_control_slave_readdata_6,
	wrclk_control_slave_readdata_7,
	altera_reset_synchronizer_int_chain_out,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_3,
	in_data_reg_0,
	in_data_reg_2,
	in_data_reg_1,
	in_data_reg_14,
	in_data_reg_8,
	in_data_reg_13,
	in_data_reg_12,
	in_data_reg_11,
	in_data_reg_10,
	in_data_reg_9,
	in_data_reg_19,
	in_data_reg_18,
	in_data_reg_17,
	in_data_reg_16,
	in_data_reg_15,
	in_data_reg_26,
	in_data_reg_21,
	in_data_reg_20,
	in_data_reg_31,
	in_data_reg_30,
	in_data_reg_29,
	in_data_reg_28,
	in_data_reg_27,
	in_data_reg_25,
	in_data_reg_24,
	in_data_reg_23,
	in_data_reg_22,
	in_data_reg_7,
	in_data_reg_6,
	in_data_reg_5,
	in_data_reg_4,
	in_data_reg_3)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARBURST_0;
input 	h2f_lw_ARBURST_1;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWID_0;
input 	h2f_lw_AWID_1;
input 	h2f_lw_AWID_2;
input 	h2f_lw_AWID_3;
input 	h2f_lw_AWID_4;
input 	h2f_lw_AWID_5;
input 	h2f_lw_AWID_6;
input 	h2f_lw_AWID_7;
input 	h2f_lw_AWID_8;
input 	h2f_lw_AWID_9;
input 	h2f_lw_AWID_10;
input 	h2f_lw_AWID_11;
input 	h2f_lw_AWLEN_0;
input 	h2f_lw_AWLEN_1;
input 	h2f_lw_AWLEN_2;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	h2f_lw_WDATA_0;
input 	h2f_lw_WDATA_1;
input 	h2f_lw_WDATA_2;
input 	h2f_lw_WDATA_3;
input 	h2f_lw_WDATA_4;
input 	h2f_lw_WDATA_5;
input 	h2f_lw_WDATA_6;
input 	h2f_lw_WDATA_7;
input 	h2f_lw_WDATA_8;
input 	h2f_lw_WDATA_9;
input 	h2f_lw_WDATA_10;
input 	h2f_lw_WDATA_11;
input 	h2f_lw_WDATA_12;
input 	h2f_lw_WDATA_13;
input 	h2f_lw_WDATA_14;
input 	h2f_lw_WDATA_15;
input 	h2f_lw_WDATA_16;
input 	h2f_lw_WDATA_17;
input 	h2f_lw_WDATA_18;
input 	h2f_lw_WDATA_19;
input 	h2f_lw_WDATA_20;
input 	h2f_lw_WDATA_21;
input 	h2f_lw_WDATA_22;
input 	h2f_lw_WDATA_23;
input 	h2f_lw_WDATA_24;
input 	h2f_lw_WDATA_25;
input 	h2f_lw_WDATA_26;
input 	h2f_lw_WDATA_27;
input 	h2f_lw_WDATA_28;
input 	h2f_lw_WDATA_29;
input 	h2f_lw_WDATA_30;
input 	h2f_lw_WDATA_31;
input 	h2f_lw_WSTRB_0;
input 	h2f_lw_WSTRB_1;
input 	h2f_lw_WSTRB_2;
input 	h2f_lw_WSTRB_3;
input 	outclk_wire_0;
output 	in_ready_hold;
output 	wait_latency_counter_0;
output 	wait_latency_counter_1;
output 	sink1_ready;
output 	ARM_A9_HPS_h2f_lw_axi_master_awready;
output 	src0_valid;
output 	source_endofpacket;
output 	src1_valid;
output 	ARM_A9_HPS_h2f_lw_axi_master_wready;
output 	mem_88_0;
output 	mem_89_0;
output 	mem_90_0;
output 	mem_91_0;
output 	mem_92_0;
output 	mem_93_0;
output 	mem_94_0;
output 	mem_95_0;
output 	mem_96_0;
output 	mem_97_0;
output 	mem_98_0;
output 	mem_99_0;
output 	out_data_0;
output 	out_data_1;
output 	out_data_2;
output 	out_data_3;
output 	out_data_4;
output 	out_data_5;
output 	out_data_6;
output 	out_data_7;
input 	r_sync_rst;
output 	m0_write;
output 	m0_read;
input 	wrclk_control_slave_readdata_0;
input 	wrclk_control_slave_readdata_1;
input 	wrclk_control_slave_readdata_2;
input 	wrclk_control_slave_readdata_3;
input 	wrclk_control_slave_readdata_4;
input 	wrclk_control_slave_readdata_5;
input 	wrclk_control_slave_readdata_6;
input 	wrclk_control_slave_readdata_7;
input 	altera_reset_synchronizer_int_chain_out;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_3;
output 	in_data_reg_0;
output 	in_data_reg_2;
output 	in_data_reg_1;
output 	in_data_reg_14;
output 	in_data_reg_8;
output 	in_data_reg_13;
output 	in_data_reg_12;
output 	in_data_reg_11;
output 	in_data_reg_10;
output 	in_data_reg_9;
output 	in_data_reg_19;
output 	in_data_reg_18;
output 	in_data_reg_17;
output 	in_data_reg_16;
output 	in_data_reg_15;
output 	in_data_reg_26;
output 	in_data_reg_21;
output 	in_data_reg_20;
output 	in_data_reg_31;
output 	in_data_reg_30;
output 	in_data_reg_29;
output 	in_data_reg_28;
output 	in_data_reg_27;
output 	in_data_reg_25;
output 	in_data_reg_24;
output 	in_data_reg_23;
output 	in_data_reg_22;
output 	in_data_reg_7;
output 	in_data_reg_6;
output 	in_data_reg_5;
output 	in_data_reg_4;
output 	in_data_reg_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arm_a9_hps_h2f_lw_axi_master_agent|Add5~1_sumout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add4~1_sumout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add5~5_sumout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add4~5_sumout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add5~9_sumout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add4~9_sumout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add5~13_sumout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add4~13_sumout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add5~17_sumout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add4~17_sumout ;
wire \cmd_mux|saved_grant[1]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem_used[1]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \fifo_hps_to_fpga_in_csr_agent|WideOr0~0_combout ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ;
wire \fifo_hps_to_fpga_in_csr_agent|cp_ready~0_combout ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \fifo_hps_to_fpga_in_csr_agent|local_write~combout ;
wire \fifo_hps_to_fpga_in_csr_agent_rsp_fifo|write~0_combout ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \cmd_mux|saved_grant[0]~q ;
wire \fifo_hps_to_fpga_in_csr_translator|read_latency_shift_reg[0]~q ;
wire \fifo_hps_to_fpga_in_csr_agent_rdata_fifo|mem_used[0]~q ;
wire \fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][112]~q ;
wire \fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem_used[0]~q ;
wire \fifo_hps_to_fpga_in_csr_agent|uncompressor|always0~0_combout ;
wire \fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][59]~q ;
wire \fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][57]~q ;
wire \fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][113]~q ;
wire \fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][69]~q ;
wire \fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][68]~q ;
wire \fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][67]~q ;
wire \fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][66]~q ;
wire \fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][65]~q ;
wire \fifo_hps_to_fpga_in_csr_agent|uncompressor|last_packet_beat~2_combout ;
wire \fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[0]~q ;
wire \fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[1]~q ;
wire \fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[2]~q ;
wire \fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[3]~q ;
wire \fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[4]~q ;
wire \fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[5]~q ;
wire \fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[6]~q ;
wire \fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[7]~q ;
wire \cmd_mux|WideOr1~combout ;
wire \cmd_mux|src_payload[0]~combout ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \fifo_hps_to_fpga_in_csr_agent|cp_ready~2_combout ;
wire \rsp_demux|WideOr0~0_combout ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ;
wire \cmd_mux|src_data[78]~combout ;
wire \cmd_mux|src_data[79]~combout ;
wire \cmd_mux|src_data[35]~combout ;
wire \cmd_mux|src_data[34]~combout ;
wire \cmd_mux|src_data[33]~combout ;
wire \cmd_mux|src_data[32]~combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|sop_enable~q ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[6]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add2~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[5]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[68]~1_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[3]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[66]~2_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[2]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[65]~3_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[4]~q ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[67]~4_combout ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[88]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[89]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ;
wire \fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ;
wire \cmd_mux|src_data[88]~combout ;
wire \cmd_mux|src_data[89]~combout ;
wire \cmd_mux|src_data[90]~combout ;
wire \cmd_mux|src_data[91]~combout ;
wire \cmd_mux|src_data[92]~combout ;
wire \cmd_mux|src_data[93]~combout ;
wire \cmd_mux|src_data[94]~combout ;
wire \cmd_mux|src_data[95]~combout ;
wire \cmd_mux|src_data[96]~combout ;
wire \cmd_mux|src_data[97]~combout ;
wire \cmd_mux|src_data[98]~combout ;
wire \cmd_mux|src_data[99]~combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[2]~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add3~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|log2ceil~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|log2ceil~1_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add1~0_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|Selector17~0_combout ;
wire \cmd_mux|src_payload~0_combout ;
wire \cmd_mux|src_data[72]~4_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[4]~1_combout ;
wire \cmd_mux|src_payload~1_combout ;
wire \cmd_mux|src_data[74]~9_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[3]~2_combout ;
wire \cmd_mux|src_data[73]~12_combout ;
wire \cmd_mux|src_payload~2_combout ;
wire \cmd_mux|src_payload~3_combout ;
wire \cmd_mux|src_payload~4_combout ;
wire \cmd_mux|src_payload~5_combout ;
wire \cmd_mux|src_payload~6_combout ;
wire \cmd_mux|src_payload~7_combout ;
wire \cmd_mux|src_payload~8_combout ;
wire \cmd_mux|src_payload~9_combout ;
wire \cmd_mux|src_payload~10_combout ;
wire \cmd_mux|src_payload~11_combout ;
wire \cmd_mux|src_payload~12_combout ;
wire \cmd_mux|src_payload~13_combout ;
wire \cmd_mux|src_payload~14_combout ;
wire \cmd_mux|src_payload~15_combout ;
wire \cmd_mux|src_payload~16_combout ;
wire \cmd_mux|src_payload~17_combout ;
wire \cmd_mux|src_payload~18_combout ;
wire \cmd_mux|src_payload~19_combout ;
wire \cmd_mux|src_payload~20_combout ;
wire \cmd_mux|src_payload~21_combout ;
wire \cmd_mux|src_payload~22_combout ;
wire \cmd_mux|src_payload~23_combout ;
wire \cmd_mux|src_payload~24_combout ;
wire \cmd_mux|src_payload~25_combout ;
wire \cmd_mux|src_payload~26_combout ;
wire \cmd_mux|src_payload~27_combout ;
wire \cmd_mux|src_payload~28_combout ;
wire \cmd_mux|src_payload~29_combout ;
wire \cmd_mux|src_payload~30_combout ;
wire \cmd_mux|src_payload~31_combout ;
wire \cmd_mux|src_payload~32_combout ;
wire \cmd_mux|src_payload~33_combout ;
wire \cmd_mux|src_data[77]~combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~3_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|Add3~1_combout ;
wire \cmd_mux|src_payload~34_combout ;
wire \cmd_mux|src_data[71]~15_combout ;
wire \arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~4_combout ;
wire \cmd_mux|src_payload~35_combout ;
wire \cmd_mux|src_data[70]~18_combout ;


Computer_System_Computer_System_mm_interconnect_1_rsp_demux rsp_demux(
	.h2f_lw_BREADY_0(h2f_lw_BREADY_0),
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.read_latency_shift_reg_0(\fifo_hps_to_fpga_in_csr_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\fifo_hps_to_fpga_in_csr_agent_rdata_fifo|mem_used[0]~q ),
	.always0(\fifo_hps_to_fpga_in_csr_agent|uncompressor|always0~0_combout ),
	.mem_59_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][57]~q ),
	.src0_valid1(src0_valid),
	.src1_valid(src1_valid),
	.WideOr0(\rsp_demux|WideOr0~0_combout ));

Computer_System_Computer_System_mm_interconnect_1_cmd_mux cmd_mux(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.h2f_lw_ARBURST_0(h2f_lw_ARBURST_0),
	.h2f_lw_ARBURST_1(h2f_lw_ARBURST_1),
	.h2f_lw_ARID_0(h2f_lw_ARID_0),
	.h2f_lw_ARID_1(h2f_lw_ARID_1),
	.h2f_lw_ARID_2(h2f_lw_ARID_2),
	.h2f_lw_ARID_3(h2f_lw_ARID_3),
	.h2f_lw_ARID_4(h2f_lw_ARID_4),
	.h2f_lw_ARID_5(h2f_lw_ARID_5),
	.h2f_lw_ARID_6(h2f_lw_ARID_6),
	.h2f_lw_ARID_7(h2f_lw_ARID_7),
	.h2f_lw_ARID_8(h2f_lw_ARID_8),
	.h2f_lw_ARID_9(h2f_lw_ARID_9),
	.h2f_lw_ARID_10(h2f_lw_ARID_10),
	.h2f_lw_ARID_11(h2f_lw_ARID_11),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWBURST_0(h2f_lw_AWBURST_0),
	.h2f_lw_AWBURST_1(h2f_lw_AWBURST_1),
	.h2f_lw_AWID_0(h2f_lw_AWID_0),
	.h2f_lw_AWID_1(h2f_lw_AWID_1),
	.h2f_lw_AWID_2(h2f_lw_AWID_2),
	.h2f_lw_AWID_3(h2f_lw_AWID_3),
	.h2f_lw_AWID_4(h2f_lw_AWID_4),
	.h2f_lw_AWID_5(h2f_lw_AWID_5),
	.h2f_lw_AWID_6(h2f_lw_AWID_6),
	.h2f_lw_AWID_7(h2f_lw_AWID_7),
	.h2f_lw_AWID_8(h2f_lw_AWID_8),
	.h2f_lw_AWID_9(h2f_lw_AWID_9),
	.h2f_lw_AWID_10(h2f_lw_AWID_10),
	.h2f_lw_AWID_11(h2f_lw_AWID_11),
	.h2f_lw_AWLEN_3(h2f_lw_AWLEN_3),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.h2f_lw_WDATA_0(h2f_lw_WDATA_0),
	.h2f_lw_WDATA_1(h2f_lw_WDATA_1),
	.h2f_lw_WDATA_2(h2f_lw_WDATA_2),
	.h2f_lw_WDATA_3(h2f_lw_WDATA_3),
	.h2f_lw_WDATA_4(h2f_lw_WDATA_4),
	.h2f_lw_WDATA_5(h2f_lw_WDATA_5),
	.h2f_lw_WDATA_6(h2f_lw_WDATA_6),
	.h2f_lw_WDATA_7(h2f_lw_WDATA_7),
	.h2f_lw_WDATA_8(h2f_lw_WDATA_8),
	.h2f_lw_WDATA_9(h2f_lw_WDATA_9),
	.h2f_lw_WDATA_10(h2f_lw_WDATA_10),
	.h2f_lw_WDATA_11(h2f_lw_WDATA_11),
	.h2f_lw_WDATA_12(h2f_lw_WDATA_12),
	.h2f_lw_WDATA_13(h2f_lw_WDATA_13),
	.h2f_lw_WDATA_14(h2f_lw_WDATA_14),
	.h2f_lw_WDATA_15(h2f_lw_WDATA_15),
	.h2f_lw_WDATA_16(h2f_lw_WDATA_16),
	.h2f_lw_WDATA_17(h2f_lw_WDATA_17),
	.h2f_lw_WDATA_18(h2f_lw_WDATA_18),
	.h2f_lw_WDATA_19(h2f_lw_WDATA_19),
	.h2f_lw_WDATA_20(h2f_lw_WDATA_20),
	.h2f_lw_WDATA_21(h2f_lw_WDATA_21),
	.h2f_lw_WDATA_22(h2f_lw_WDATA_22),
	.h2f_lw_WDATA_23(h2f_lw_WDATA_23),
	.h2f_lw_WDATA_24(h2f_lw_WDATA_24),
	.h2f_lw_WDATA_25(h2f_lw_WDATA_25),
	.h2f_lw_WDATA_26(h2f_lw_WDATA_26),
	.h2f_lw_WDATA_27(h2f_lw_WDATA_27),
	.h2f_lw_WDATA_28(h2f_lw_WDATA_28),
	.h2f_lw_WDATA_29(h2f_lw_WDATA_29),
	.h2f_lw_WDATA_30(h2f_lw_WDATA_30),
	.h2f_lw_WDATA_31(h2f_lw_WDATA_31),
	.h2f_lw_WSTRB_0(h2f_lw_WSTRB_0),
	.h2f_lw_WSTRB_1(h2f_lw_WSTRB_1),
	.h2f_lw_WSTRB_2(h2f_lw_WSTRB_2),
	.h2f_lw_WSTRB_3(h2f_lw_WSTRB_3),
	.outclk_wire_0(outclk_wire_0),
	.Add5(\arm_a9_hps_h2f_lw_axi_master_agent|Add5~1_sumout ),
	.Add4(\arm_a9_hps_h2f_lw_axi_master_agent|Add4~1_sumout ),
	.Add51(\arm_a9_hps_h2f_lw_axi_master_agent|Add5~5_sumout ),
	.Add41(\arm_a9_hps_h2f_lw_axi_master_agent|Add4~5_sumout ),
	.Add52(\arm_a9_hps_h2f_lw_axi_master_agent|Add5~9_sumout ),
	.Add42(\arm_a9_hps_h2f_lw_axi_master_agent|Add4~9_sumout ),
	.Add53(\arm_a9_hps_h2f_lw_axi_master_agent|Add5~13_sumout ),
	.Add43(\arm_a9_hps_h2f_lw_axi_master_agent|Add4~13_sumout ),
	.Add54(\arm_a9_hps_h2f_lw_axi_master_agent|Add5~17_sumout ),
	.Add44(\arm_a9_hps_h2f_lw_axi_master_agent|Add4~17_sumout ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.nxt_in_ready(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready1(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.sink1_ready1(sink1_ready),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.r_sync_rst(r_sync_rst),
	.WideOr11(\cmd_mux|WideOr1~combout ),
	.src_payload_0(\cmd_mux|src_payload[0]~combout ),
	.src_data_78(\cmd_mux|src_data[78]~combout ),
	.src_data_79(\cmd_mux|src_data[79]~combout ),
	.src_data_35(\cmd_mux|src_data[35]~combout ),
	.src_data_34(\cmd_mux|src_data[34]~combout ),
	.src_data_33(\cmd_mux|src_data[33]~combout ),
	.src_data_32(\cmd_mux|src_data[32]~combout ),
	.src_data_88(\cmd_mux|src_data[88]~combout ),
	.src_data_89(\cmd_mux|src_data[89]~combout ),
	.src_data_90(\cmd_mux|src_data[90]~combout ),
	.src_data_91(\cmd_mux|src_data[91]~combout ),
	.src_data_92(\cmd_mux|src_data[92]~combout ),
	.src_data_93(\cmd_mux|src_data[93]~combout ),
	.src_data_94(\cmd_mux|src_data[94]~combout ),
	.src_data_95(\cmd_mux|src_data[95]~combout ),
	.src_data_96(\cmd_mux|src_data[96]~combout ),
	.src_data_97(\cmd_mux|src_data[97]~combout ),
	.src_data_98(\cmd_mux|src_data[98]~combout ),
	.src_data_99(\cmd_mux|src_data[99]~combout ),
	.Add3(\arm_a9_hps_h2f_lw_axi_master_agent|Add3~0_combout ),
	.log2ceil(\arm_a9_hps_h2f_lw_axi_master_agent|log2ceil~0_combout ),
	.log2ceil1(\arm_a9_hps_h2f_lw_axi_master_agent|log2ceil~1_combout ),
	.Add1(\arm_a9_hps_h2f_lw_axi_master_agent|Add1~0_combout ),
	.Selector17(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|Selector17~0_combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.src_data_72(\cmd_mux|src_data[72]~4_combout ),
	.src_payload1(\cmd_mux|src_payload~1_combout ),
	.src_data_74(\cmd_mux|src_data[74]~9_combout ),
	.src_data_73(\cmd_mux|src_data[73]~12_combout ),
	.src_payload2(\cmd_mux|src_payload~2_combout ),
	.src_payload3(\cmd_mux|src_payload~3_combout ),
	.src_payload4(\cmd_mux|src_payload~4_combout ),
	.src_payload5(\cmd_mux|src_payload~5_combout ),
	.src_payload6(\cmd_mux|src_payload~6_combout ),
	.src_payload7(\cmd_mux|src_payload~7_combout ),
	.src_payload8(\cmd_mux|src_payload~8_combout ),
	.src_payload9(\cmd_mux|src_payload~9_combout ),
	.src_payload10(\cmd_mux|src_payload~10_combout ),
	.src_payload11(\cmd_mux|src_payload~11_combout ),
	.src_payload12(\cmd_mux|src_payload~12_combout ),
	.src_payload13(\cmd_mux|src_payload~13_combout ),
	.src_payload14(\cmd_mux|src_payload~14_combout ),
	.src_payload15(\cmd_mux|src_payload~15_combout ),
	.src_payload16(\cmd_mux|src_payload~16_combout ),
	.src_payload17(\cmd_mux|src_payload~17_combout ),
	.src_payload18(\cmd_mux|src_payload~18_combout ),
	.src_payload19(\cmd_mux|src_payload~19_combout ),
	.src_payload20(\cmd_mux|src_payload~20_combout ),
	.src_payload21(\cmd_mux|src_payload~21_combout ),
	.src_payload22(\cmd_mux|src_payload~22_combout ),
	.src_payload23(\cmd_mux|src_payload~23_combout ),
	.src_payload24(\cmd_mux|src_payload~24_combout ),
	.src_payload25(\cmd_mux|src_payload~25_combout ),
	.src_payload26(\cmd_mux|src_payload~26_combout ),
	.src_payload27(\cmd_mux|src_payload~27_combout ),
	.src_payload28(\cmd_mux|src_payload~28_combout ),
	.src_payload29(\cmd_mux|src_payload~29_combout ),
	.src_payload30(\cmd_mux|src_payload~30_combout ),
	.src_payload31(\cmd_mux|src_payload~31_combout ),
	.src_payload32(\cmd_mux|src_payload~32_combout ),
	.src_payload33(\cmd_mux|src_payload~33_combout ),
	.src_data_77(\cmd_mux|src_data[77]~combout ),
	.Add31(\arm_a9_hps_h2f_lw_axi_master_agent|Add3~1_combout ),
	.src_payload34(\cmd_mux|src_payload~34_combout ),
	.src_data_71(\cmd_mux|src_data[71]~15_combout ),
	.src_payload35(\cmd_mux|src_payload~35_combout ),
	.src_data_70(\cmd_mux|src_data[70]~18_combout ));

Computer_System_altera_merlin_burst_adapter_2 fifo_hps_to_fpga_in_csr_burst_adapter(
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARADDR_4(h2f_lw_ARADDR_4),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.outclk_wire_0(outclk_wire_0),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.stateST_COMP_TRANS(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.in_ready_hold(in_ready_hold),
	.stateST_UNCOMP_WR_SUBBURST(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.out_valid_reg(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\fifo_hps_to_fpga_in_csr_agent|WideOr0~0_combout ),
	.wait_latency_counter_0(wait_latency_counter_0),
	.in_data_reg_59(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.cp_ready(\fifo_hps_to_fpga_in_csr_agent|cp_ready~0_combout ),
	.nxt_in_ready(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.local_write(\fifo_hps_to_fpga_in_csr_agent|local_write~combout ),
	.write(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|write~0_combout ),
	.nxt_in_ready1(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.r_sync_rst(r_sync_rst),
	.WideOr1(\cmd_mux|WideOr1~combout ),
	.src_payload_0(\cmd_mux|src_payload[0]~combout ),
	.nxt_out_eop(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_uncomp_byte_cnt_reg_5(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_byte_cnt_reg_2(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.cp_ready1(\fifo_hps_to_fpga_in_csr_agent|cp_ready~2_combout ),
	.in_data_reg_60(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.src_data_78(\cmd_mux|src_data[78]~combout ),
	.src_data_79(\cmd_mux|src_data[79]~combout ),
	.src_data_35(\cmd_mux|src_data[35]~combout ),
	.src_data_34(\cmd_mux|src_data[34]~combout ),
	.src_data_33(\cmd_mux|src_data[33]~combout ),
	.src_data_32(\cmd_mux|src_data[32]~combout ),
	.sop_enable(\arm_a9_hps_h2f_lw_axi_master_agent|sop_enable~q ),
	.burst_bytecount_6(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[6]~q ),
	.write_cp_data_69(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ),
	.Add2(\arm_a9_hps_h2f_lw_axi_master_agent|Add2~0_combout ),
	.burst_bytecount_5(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[5]~q ),
	.write_cp_data_68(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[68]~1_combout ),
	.burst_bytecount_3(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[3]~q ),
	.write_cp_data_66(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[66]~2_combout ),
	.burst_bytecount_2(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[2]~q ),
	.write_cp_data_65(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[65]~3_combout ),
	.burst_bytecount_4(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[4]~q ),
	.write_cp_data_67(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[67]~4_combout ),
	.in_data_reg_88(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[88]~q ),
	.in_data_reg_89(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[89]~q ),
	.in_data_reg_90(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ),
	.in_data_reg_91(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.in_data_reg_92(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.src_data_88(\cmd_mux|src_data[88]~combout ),
	.src_data_89(\cmd_mux|src_data[89]~combout ),
	.src_data_90(\cmd_mux|src_data[90]~combout ),
	.src_data_91(\cmd_mux|src_data[91]~combout ),
	.src_data_92(\cmd_mux|src_data[92]~combout ),
	.src_data_93(\cmd_mux|src_data[93]~combout ),
	.src_data_94(\cmd_mux|src_data[94]~combout ),
	.src_data_95(\cmd_mux|src_data[95]~combout ),
	.src_data_96(\cmd_mux|src_data[96]~combout ),
	.src_data_97(\cmd_mux|src_data[97]~combout ),
	.src_data_98(\cmd_mux|src_data[98]~combout ),
	.src_data_99(\cmd_mux|src_data[99]~combout ),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_4(int_nxt_addr_reg_dly_4),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.out_data_2(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[2]~0_combout ),
	.src_data_72(\cmd_mux|src_data[72]~4_combout ),
	.out_data_4(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[4]~1_combout ),
	.src_data_74(\cmd_mux|src_data[74]~9_combout ),
	.out_data_3(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[3]~2_combout ),
	.src_data_73(\cmd_mux|src_data[73]~12_combout ),
	.in_data_reg_0(in_data_reg_0),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_31(in_data_reg_31),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_24(in_data_reg_24),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_3(in_data_reg_3),
	.src_payload(\cmd_mux|src_payload~2_combout ),
	.src_payload1(\cmd_mux|src_payload~3_combout ),
	.src_payload2(\cmd_mux|src_payload~4_combout ),
	.src_payload3(\cmd_mux|src_payload~5_combout ),
	.src_payload4(\cmd_mux|src_payload~6_combout ),
	.src_payload5(\cmd_mux|src_payload~7_combout ),
	.src_payload6(\cmd_mux|src_payload~8_combout ),
	.src_payload7(\cmd_mux|src_payload~9_combout ),
	.src_payload8(\cmd_mux|src_payload~10_combout ),
	.src_payload9(\cmd_mux|src_payload~11_combout ),
	.src_payload10(\cmd_mux|src_payload~12_combout ),
	.src_payload11(\cmd_mux|src_payload~13_combout ),
	.src_payload12(\cmd_mux|src_payload~14_combout ),
	.src_payload13(\cmd_mux|src_payload~15_combout ),
	.src_payload14(\cmd_mux|src_payload~16_combout ),
	.src_payload15(\cmd_mux|src_payload~17_combout ),
	.src_payload16(\cmd_mux|src_payload~18_combout ),
	.src_payload17(\cmd_mux|src_payload~19_combout ),
	.src_payload18(\cmd_mux|src_payload~20_combout ),
	.src_payload19(\cmd_mux|src_payload~21_combout ),
	.src_payload20(\cmd_mux|src_payload~22_combout ),
	.src_payload21(\cmd_mux|src_payload~23_combout ),
	.src_payload22(\cmd_mux|src_payload~24_combout ),
	.src_payload23(\cmd_mux|src_payload~25_combout ),
	.src_payload24(\cmd_mux|src_payload~26_combout ),
	.src_payload25(\cmd_mux|src_payload~27_combout ),
	.src_payload26(\cmd_mux|src_payload~28_combout ),
	.src_payload27(\cmd_mux|src_payload~29_combout ),
	.src_payload28(\cmd_mux|src_payload~30_combout ),
	.src_payload29(\cmd_mux|src_payload~31_combout ),
	.src_payload30(\cmd_mux|src_payload~32_combout ),
	.src_payload31(\cmd_mux|src_payload~33_combout ),
	.src_data_77(\cmd_mux|src_data[77]~combout ),
	.out_data_1(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~3_combout ),
	.src_data_71(\cmd_mux|src_data[71]~15_combout ),
	.out_data_0(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~4_combout ),
	.src_data_70(\cmd_mux|src_data[70]~18_combout ));

Computer_System_altera_avalon_sc_fifo_4 fifo_hps_to_fpga_in_csr_agent_rdata_fifo(
	.clk(outclk_wire_0),
	.read_latency_shift_reg_0(\fifo_hps_to_fpga_in_csr_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\fifo_hps_to_fpga_in_csr_agent_rdata_fifo|mem_used[0]~q ),
	.mem_112_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_01(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[0]~q ),
	.out_data_0(out_data_0),
	.av_readdata_pre_1(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[1]~q ),
	.out_data_1(out_data_1),
	.av_readdata_pre_2(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[2]~q ),
	.out_data_2(out_data_2),
	.av_readdata_pre_3(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[3]~q ),
	.out_data_3(out_data_3),
	.av_readdata_pre_4(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[4]~q ),
	.out_data_4(out_data_4),
	.av_readdata_pre_5(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[5]~q ),
	.out_data_5(out_data_5),
	.av_readdata_pre_6(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[6]~q ),
	.out_data_6(out_data_6),
	.av_readdata_pre_7(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[7]~q ),
	.out_data_7(out_data_7),
	.reset(r_sync_rst),
	.WideOr0(\rsp_demux|WideOr0~0_combout ));

Computer_System_altera_avalon_sc_fifo_5 fifo_hps_to_fpga_in_csr_agent_rsp_fifo(
	.clk(outclk_wire_0),
	.stateST_UNCOMP_WR_SUBBURST(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.out_valid_reg(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\fifo_hps_to_fpga_in_csr_agent|WideOr0~0_combout ),
	.wait_latency_counter_0(wait_latency_counter_0),
	.in_data_reg_59(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.cp_ready(\fifo_hps_to_fpga_in_csr_agent|cp_ready~0_combout ),
	.local_write(\fifo_hps_to_fpga_in_csr_agent|local_write~combout ),
	.write(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|write~0_combout ),
	.read_latency_shift_reg_0(\fifo_hps_to_fpga_in_csr_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\fifo_hps_to_fpga_in_csr_agent_rdata_fifo|mem_used[0]~q ),
	.mem_112_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_01(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem_used[0]~q ),
	.mem_59_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][57]~q ),
	.mem_113_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][113]~q ),
	.mem_69_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat(\fifo_hps_to_fpga_in_csr_agent|uncompressor|last_packet_beat~2_combout ),
	.mem_88_0(mem_88_0),
	.mem_89_0(mem_89_0),
	.mem_90_0(mem_90_0),
	.mem_91_0(mem_91_0),
	.mem_92_0(mem_92_0),
	.mem_93_0(mem_93_0),
	.mem_94_0(mem_94_0),
	.mem_95_0(mem_95_0),
	.mem_96_0(mem_96_0),
	.mem_97_0(mem_97_0),
	.mem_98_0(mem_98_0),
	.mem_99_0(mem_99_0),
	.reset(r_sync_rst),
	.nxt_out_eop(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.out_uncomp_byte_cnt_reg_5(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_byte_cnt_reg_2(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.WideOr01(\rsp_demux|WideOr0~0_combout ),
	.in_data_reg_60(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.in_data_reg_88(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[88]~q ),
	.in_data_reg_89(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[89]~q ),
	.in_data_reg_90(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[90]~q ),
	.in_data_reg_91(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[91]~q ),
	.in_data_reg_92(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ));

Computer_System_altera_merlin_slave_agent_2 fifo_hps_to_fpga_in_csr_agent(
	.outclk_wire_0(outclk_wire_0),
	.stateST_COMP_TRANS(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.in_ready_hold(in_ready_hold),
	.out_valid_reg(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\fifo_hps_to_fpga_in_csr_agent|WideOr0~0_combout ),
	.wait_latency_counter_0(wait_latency_counter_0),
	.in_data_reg_59(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.wait_latency_counter_1(wait_latency_counter_1),
	.cp_ready(\fifo_hps_to_fpga_in_csr_agent|cp_ready~0_combout ),
	.local_write1(\fifo_hps_to_fpga_in_csr_agent|local_write~combout ),
	.read_latency_shift_reg_0(\fifo_hps_to_fpga_in_csr_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\fifo_hps_to_fpga_in_csr_agent_rdata_fifo|mem_used[0]~q ),
	.mem_112_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][112]~q ),
	.mem_used_01(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem_used[0]~q ),
	.always0(\fifo_hps_to_fpga_in_csr_agent|uncompressor|always0~0_combout ),
	.mem_57_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][57]~q ),
	.mem_113_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][113]~q ),
	.mem_69_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\fifo_hps_to_fpga_in_csr_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat(\fifo_hps_to_fpga_in_csr_agent|uncompressor|last_packet_beat~2_combout ),
	.source_endofpacket(source_endofpacket),
	.r_sync_rst(r_sync_rst),
	.cp_ready1(\fifo_hps_to_fpga_in_csr_agent|cp_ready~2_combout ),
	.WideOr01(\rsp_demux|WideOr0~0_combout ),
	.in_data_reg_60(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.m0_write1(m0_write),
	.m0_read(m0_read));

Computer_System_altera_merlin_axi_master_ni_1 arm_a9_hps_h2f_lw_axi_master_agent(
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWADDR_0(h2f_lw_AWADDR_0),
	.h2f_lw_AWADDR_1(h2f_lw_AWADDR_1),
	.h2f_lw_AWADDR_2(h2f_lw_AWADDR_2),
	.h2f_lw_AWADDR_3(h2f_lw_AWADDR_3),
	.h2f_lw_AWADDR_4(h2f_lw_AWADDR_4),
	.h2f_lw_AWBURST_0(h2f_lw_AWBURST_0),
	.h2f_lw_AWBURST_1(h2f_lw_AWBURST_1),
	.h2f_lw_AWLEN_0(h2f_lw_AWLEN_0),
	.h2f_lw_AWLEN_1(h2f_lw_AWLEN_1),
	.h2f_lw_AWLEN_2(h2f_lw_AWLEN_2),
	.h2f_lw_AWLEN_3(h2f_lw_AWLEN_3),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.outclk_wire_0(outclk_wire_0),
	.Add5(\arm_a9_hps_h2f_lw_axi_master_agent|Add5~1_sumout ),
	.Add4(\arm_a9_hps_h2f_lw_axi_master_agent|Add4~1_sumout ),
	.Add51(\arm_a9_hps_h2f_lw_axi_master_agent|Add5~5_sumout ),
	.Add41(\arm_a9_hps_h2f_lw_axi_master_agent|Add4~5_sumout ),
	.Add52(\arm_a9_hps_h2f_lw_axi_master_agent|Add5~9_sumout ),
	.Add42(\arm_a9_hps_h2f_lw_axi_master_agent|Add4~9_sumout ),
	.Add53(\arm_a9_hps_h2f_lw_axi_master_agent|Add5~13_sumout ),
	.Add43(\arm_a9_hps_h2f_lw_axi_master_agent|Add4~13_sumout ),
	.Add54(\arm_a9_hps_h2f_lw_axi_master_agent|Add5~17_sumout ),
	.Add44(\arm_a9_hps_h2f_lw_axi_master_agent|Add4~17_sumout ),
	.nxt_in_ready(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready1(\fifo_hps_to_fpga_in_csr_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_0(\cmd_mux|saved_grant[0]~q ),
	.awready(ARM_A9_HPS_h2f_lw_axi_master_awready),
	.wready(ARM_A9_HPS_h2f_lw_axi_master_wready),
	.sop_enable1(\arm_a9_hps_h2f_lw_axi_master_agent|sop_enable~q ),
	.burst_bytecount_6(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[6]~q ),
	.write_cp_data_69(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ),
	.Add2(\arm_a9_hps_h2f_lw_axi_master_agent|Add2~0_combout ),
	.burst_bytecount_5(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[5]~q ),
	.write_cp_data_68(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[68]~1_combout ),
	.burst_bytecount_3(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[3]~q ),
	.write_cp_data_66(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[66]~2_combout ),
	.burst_bytecount_2(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[2]~q ),
	.write_cp_data_65(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[65]~3_combout ),
	.burst_bytecount_4(\arm_a9_hps_h2f_lw_axi_master_agent|burst_bytecount[4]~q ),
	.write_cp_data_67(\arm_a9_hps_h2f_lw_axi_master_agent|write_cp_data[67]~4_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.out_data_2(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[2]~0_combout ),
	.Add3(\arm_a9_hps_h2f_lw_axi_master_agent|Add3~0_combout ),
	.log2ceil(\arm_a9_hps_h2f_lw_axi_master_agent|log2ceil~0_combout ),
	.log2ceil1(\arm_a9_hps_h2f_lw_axi_master_agent|log2ceil~1_combout ),
	.Add1(\arm_a9_hps_h2f_lw_axi_master_agent|Add1~0_combout ),
	.Selector17(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|Selector17~0_combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.out_data_4(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[4]~1_combout ),
	.src_payload1(\cmd_mux|src_payload~1_combout ),
	.out_data_3(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[3]~2_combout ),
	.out_data_1(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~3_combout ),
	.Add31(\arm_a9_hps_h2f_lw_axi_master_agent|Add3~1_combout ),
	.src_payload2(\cmd_mux|src_payload~34_combout ),
	.out_data_0(\arm_a9_hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~4_combout ),
	.src_payload3(\cmd_mux|src_payload~35_combout ));

Computer_System_altera_merlin_slave_translator_2 fifo_hps_to_fpga_in_csr_translator(
	.clk(outclk_wire_0),
	.in_ready_hold(in_ready_hold),
	.wait_latency_counter_0(wait_latency_counter_0),
	.wait_latency_counter_1(wait_latency_counter_1),
	.cp_ready(\fifo_hps_to_fpga_in_csr_agent|cp_ready~0_combout ),
	.read_latency_shift_reg_0(\fifo_hps_to_fpga_in_csr_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\fifo_hps_to_fpga_in_csr_translator|av_readdata_pre[7]~q ),
	.reset(r_sync_rst),
	.m0_write(m0_write),
	.m0_read(m0_read),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,wrclk_control_slave_readdata_7,wrclk_control_slave_readdata_6,wrclk_control_slave_readdata_5,wrclk_control_slave_readdata_4,wrclk_control_slave_readdata_3,wrclk_control_slave_readdata_2,
wrclk_control_slave_readdata_1,wrclk_control_slave_readdata_0}));

endmodule

module Computer_System_altera_avalon_sc_fifo_4 (
	clk,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_112_0,
	mem_used_01,
	av_readdata_pre_0,
	out_data_0,
	av_readdata_pre_1,
	out_data_1,
	av_readdata_pre_2,
	out_data_2,
	av_readdata_pre_3,
	out_data_3,
	av_readdata_pre_4,
	out_data_4,
	av_readdata_pre_5,
	out_data_5,
	av_readdata_pre_6,
	out_data_6,
	av_readdata_pre_7,
	out_data_7,
	reset,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_112_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	out_data_0;
input 	av_readdata_pre_1;
output 	out_data_1;
input 	av_readdata_pre_2;
output 	out_data_2;
input 	av_readdata_pre_3;
output 	out_data_3;
input 	av_readdata_pre_4;
output 	out_data_4;
input 	av_readdata_pre_5;
output 	out_data_5;
input 	av_readdata_pre_6;
output 	out_data_6;
input 	av_readdata_pre_7;
output 	out_data_7;
input 	reset;
input 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[0][0]~q ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[0][1]~q ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[0][2]~q ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[0][3]~q ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[0][4]~q ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[0][5]~q ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[0][6]~q ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[0][7]~q ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \out_data[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_0),
	.datad(!\mem[0][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[0]~0 .extended_lut = "off";
defparam \out_data[0]~0 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \out_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_1),
	.datad(!\mem[0][1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[1]~1 .extended_lut = "off";
defparam \out_data[1]~1 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \out_data[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[2]~2 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_2),
	.datad(!\mem[0][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[2]~2 .extended_lut = "off";
defparam \out_data[2]~2 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \out_data[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \out_data[3]~3 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_3),
	.datad(!\mem[0][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[3]~3 .extended_lut = "off";
defparam \out_data[3]~3 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \out_data[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \out_data[4]~4 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_4),
	.datad(!\mem[0][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[4]~4 .extended_lut = "off";
defparam \out_data[4]~4 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \out_data[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \out_data[5]~5 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_5),
	.datad(!\mem[0][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[5]~5 .extended_lut = "off";
defparam \out_data[5]~5 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \out_data[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \out_data[6]~6 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_6),
	.datad(!\mem[0][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[6]~6 .extended_lut = "off";
defparam \out_data[6]~6 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \out_data[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \out_data[7]~7 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!av_readdata_pre_7),
	.datad(!\mem[0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[7]~7 .extended_lut = "off";
defparam \out_data[7]~7 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \out_data[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][0]~q ),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][1]~q ),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][2]~q ),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][3]~q ),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][4]~q ),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][5]~q ),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][6]~q ),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!av_readdata_pre_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\mem[0][7]~q ),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

endmodule

module Computer_System_altera_avalon_sc_fifo_5 (
	clk,
	stateST_UNCOMP_WR_SUBBURST,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_0,
	in_data_reg_59,
	cp_ready,
	local_write,
	write,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_112_0,
	mem_used_01,
	mem_59_0,
	mem_57_0,
	mem_113_0,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat,
	mem_88_0,
	mem_89_0,
	mem_90_0,
	mem_91_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	reset,
	nxt_out_eop,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	WideOr01,
	in_data_reg_60,
	in_data_reg_88,
	in_data_reg_89,
	in_data_reg_90,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	stateST_UNCOMP_WR_SUBBURST;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	wait_latency_counter_0;
input 	in_data_reg_59;
input 	cp_ready;
input 	local_write;
output 	write;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
output 	mem_112_0;
output 	mem_used_01;
output 	mem_59_0;
output 	mem_57_0;
output 	mem_113_0;
output 	mem_69_0;
output 	mem_68_0;
output 	mem_67_0;
output 	mem_66_0;
output 	mem_65_0;
input 	last_packet_beat;
output 	mem_88_0;
output 	mem_89_0;
output 	mem_90_0;
output 	mem_91_0;
output 	mem_92_0;
output 	mem_93_0;
output 	mem_94_0;
output 	mem_95_0;
output 	mem_96_0;
output 	mem_97_0;
output 	mem_98_0;
output 	mem_99_0;
input 	reset;
input 	nxt_out_eop;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_6;
input 	WideOr01;
input 	in_data_reg_60;
input 	in_data_reg_88;
input 	in_data_reg_89;
input 	in_data_reg_90;
input 	in_data_reg_91;
input 	in_data_reg_92;
input 	in_data_reg_93;
input 	in_data_reg_94;
input 	in_data_reg_95;
input 	in_data_reg_96;
input 	in_data_reg_97;
input 	in_data_reg_98;
input 	in_data_reg_99;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \write~1_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][112]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][59]~q ;
wire \mem~0_combout ;
wire \mem[1][60]~q ;
wire \mem~1_combout ;
wire \mem[1][113]~q ;
wire \mem~2_combout ;
wire \mem[1][69]~q ;
wire \mem~3_combout ;
wire \mem[1][68]~q ;
wire \mem~4_combout ;
wire \mem[1][67]~q ;
wire \mem~5_combout ;
wire \mem[1][66]~q ;
wire \mem~6_combout ;
wire \mem[1][65]~q ;
wire \mem~7_combout ;
wire \mem[1][88]~q ;
wire \mem~8_combout ;
wire \mem[1][89]~q ;
wire \mem~9_combout ;
wire \mem[1][90]~q ;
wire \mem~10_combout ;
wire \mem[1][91]~q ;
wire \mem~11_combout ;
wire \mem[1][92]~q ;
wire \mem~12_combout ;
wire \mem[1][93]~q ;
wire \mem~13_combout ;
wire \mem[1][94]~q ;
wire \mem~14_combout ;
wire \mem[1][95]~q ;
wire \mem~15_combout ;
wire \mem[1][96]~q ;
wire \mem~16_combout ;
wire \mem[1][97]~q ;
wire \mem~17_combout ;
wire \mem[1][98]~q ;
wire \mem~18_combout ;
wire \mem[1][99]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!wait_latency_counter_0),
	.datad(!local_write),
	.datae(!cp_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h88888AA888888AA8;
defparam \write~0 .shared_arith = "off";

dffeas \mem[0][112] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_112_0),
	.prn(vcc));
defparam \mem[0][112] .is_wysiwyg = "true";
defparam \mem[0][112] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_01),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][59] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_59_0),
	.prn(vcc));
defparam \mem[0][59] .is_wysiwyg = "true";
defparam \mem[0][59] .power_up = "low";

dffeas \mem[0][57] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_57_0),
	.prn(vcc));
defparam \mem[0][57] .is_wysiwyg = "true";
defparam \mem[0][57] .power_up = "low";

dffeas \mem[0][113] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_113_0),
	.prn(vcc));
defparam \mem[0][113] .is_wysiwyg = "true";
defparam \mem[0][113] .power_up = "low";

dffeas \mem[0][69] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_69_0),
	.prn(vcc));
defparam \mem[0][69] .is_wysiwyg = "true";
defparam \mem[0][69] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][65] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_65_0),
	.prn(vcc));
defparam \mem[0][65] .is_wysiwyg = "true";
defparam \mem[0][65] .power_up = "low";

dffeas \mem[0][88] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_88_0),
	.prn(vcc));
defparam \mem[0][88] .is_wysiwyg = "true";
defparam \mem[0][88] .power_up = "low";

dffeas \mem[0][89] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_89_0),
	.prn(vcc));
defparam \mem[0][89] .is_wysiwyg = "true";
defparam \mem[0][89] .power_up = "low";

dffeas \mem[0][90] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_90_0),
	.prn(vcc));
defparam \mem[0][90] .is_wysiwyg = "true";
defparam \mem[0][90] .power_up = "low";

dffeas \mem[0][91] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_91_0),
	.prn(vcc));
defparam \mem[0][91] .is_wysiwyg = "true";
defparam \mem[0][91] .power_up = "low";

dffeas \mem[0][92] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_92_0),
	.prn(vcc));
defparam \mem[0][92] .is_wysiwyg = "true";
defparam \mem[0][92] .power_up = "low";

dffeas \mem[0][93] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_93_0),
	.prn(vcc));
defparam \mem[0][93] .is_wysiwyg = "true";
defparam \mem[0][93] .power_up = "low";

dffeas \mem[0][94] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_94_0),
	.prn(vcc));
defparam \mem[0][94] .is_wysiwyg = "true";
defparam \mem[0][94] .power_up = "low";

dffeas \mem[0][95] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_95_0),
	.prn(vcc));
defparam \mem[0][95] .is_wysiwyg = "true";
defparam \mem[0][95] .power_up = "low";

dffeas \mem[0][96] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_96_0),
	.prn(vcc));
defparam \mem[0][96] .is_wysiwyg = "true";
defparam \mem[0][96] .power_up = "low";

dffeas \mem[0][97] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_97_0),
	.prn(vcc));
defparam \mem[0][97] .is_wysiwyg = "true";
defparam \mem[0][97] .power_up = "low";

dffeas \mem[0][98] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_98_0),
	.prn(vcc));
defparam \mem[0][98] .is_wysiwyg = "true";
defparam \mem[0][98] .power_up = "low";

dffeas \mem[0][99] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_99_0),
	.prn(vcc));
defparam \mem[0][99] .is_wysiwyg = "true";
defparam \mem[0][99] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!last_packet_beat),
	.datae(!WideOr01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h00007F0000007F00;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!out_valid_reg),
	.datab(!in_data_reg_59),
	.datac(!write),
	.datad(!nxt_out_eop),
	.datae(!in_data_reg_60),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0001050500010505;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_01),
	.datac(!\read~0_combout ),
	.datad(!\write~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5431543154315431;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][112] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][112]~q ),
	.prn(vcc));
defparam \mem[1][112] .is_wysiwyg = "true";
defparam \mem[1][112] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!in_data_reg_59),
	.datac(!\mem[1][112]~q ),
	.datad(!out_valid_reg),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_60),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h000A0F0F003B0F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_01),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_01),
	.datac(!\read~0_combout ),
	.datad(!\write~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h31FF31FF31FF31FF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][59] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][59]~q ),
	.prn(vcc));
defparam \mem[1][59] .is_wysiwyg = "true";
defparam \mem[1][59] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_59),
	.datac(!\mem[1][59]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][60] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][60]~q ),
	.prn(vcc));
defparam \mem[1][60] .is_wysiwyg = "true";
defparam \mem[1][60] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_60),
	.datac(!\mem[1][60]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][113] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][113]~q ),
	.prn(vcc));
defparam \mem[1][113] .is_wysiwyg = "true";
defparam \mem[1][113] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][113]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][69]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0437043704370437;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][68]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0437043704370437;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][67]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0437043704370437;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0437043704370437;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][65] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][65]~q ),
	.prn(vcc));
defparam \mem[1][65] .is_wysiwyg = "true";
defparam \mem[1][65] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!stateST_UNCOMP_WR_SUBBURST),
	.datab(!mem_used_1),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\mem[1][65]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h048C37BF048C37BF;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][88] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][88]~q ),
	.prn(vcc));
defparam \mem[1][88] .is_wysiwyg = "true";
defparam \mem[1][88] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][88]~q ),
	.datac(!in_data_reg_88),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][89] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][89]~q ),
	.prn(vcc));
defparam \mem[1][89] .is_wysiwyg = "true";
defparam \mem[1][89] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][89]~q ),
	.datac(!in_data_reg_89),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][90] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][90]~q ),
	.prn(vcc));
defparam \mem[1][90] .is_wysiwyg = "true";
defparam \mem[1][90] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][90]~q ),
	.datac(!in_data_reg_90),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][91] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][91]~q ),
	.prn(vcc));
defparam \mem[1][91] .is_wysiwyg = "true";
defparam \mem[1][91] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][91]~q ),
	.datac(!in_data_reg_91),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][92] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][92]~q ),
	.prn(vcc));
defparam \mem[1][92] .is_wysiwyg = "true";
defparam \mem[1][92] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][92]~q ),
	.datac(!in_data_reg_92),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][93] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][93]~q ),
	.prn(vcc));
defparam \mem[1][93] .is_wysiwyg = "true";
defparam \mem[1][93] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][93]~q ),
	.datac(!in_data_reg_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(!in_data_reg_94),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][95] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][95]~q ),
	.prn(vcc));
defparam \mem[1][95] .is_wysiwyg = "true";
defparam \mem[1][95] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][95]~q ),
	.datac(!in_data_reg_95),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][96] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][96]~q ),
	.prn(vcc));
defparam \mem[1][96] .is_wysiwyg = "true";
defparam \mem[1][96] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][96]~q ),
	.datac(!in_data_reg_96),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][97] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][97]~q ),
	.prn(vcc));
defparam \mem[1][97] .is_wysiwyg = "true";
defparam \mem[1][97] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][97]~q ),
	.datac(!in_data_reg_97),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][98] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][98]~q ),
	.prn(vcc));
defparam \mem[1][98] .is_wysiwyg = "true";
defparam \mem[1][98] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][98]~q ),
	.datac(!in_data_reg_98),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][99] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][99]~q ),
	.prn(vcc));
defparam \mem[1][99] .is_wysiwyg = "true";
defparam \mem[1][99] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][99]~q ),
	.datac(!in_data_reg_99),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_axi_master_ni_1 (
	h2f_lw_AWVALID_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	outclk_wire_0,
	Add5,
	Add4,
	Add51,
	Add41,
	Add52,
	Add42,
	Add53,
	Add43,
	Add54,
	Add44,
	nxt_in_ready,
	nxt_in_ready1,
	saved_grant_0,
	awready,
	wready,
	sop_enable1,
	burst_bytecount_6,
	write_cp_data_69,
	Add2,
	burst_bytecount_5,
	write_cp_data_68,
	burst_bytecount_3,
	write_cp_data_66,
	burst_bytecount_2,
	write_cp_data_65,
	burst_bytecount_4,
	write_cp_data_67,
	altera_reset_synchronizer_int_chain_out,
	out_data_2,
	Add3,
	log2ceil,
	log2ceil1,
	Add1,
	Selector17,
	src_payload,
	out_data_4,
	src_payload1,
	out_data_3,
	out_data_1,
	Add31,
	src_payload2,
	out_data_0,
	src_payload3)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWLEN_0;
input 	h2f_lw_AWLEN_1;
input 	h2f_lw_AWLEN_2;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	outclk_wire_0;
output 	Add5;
output 	Add4;
output 	Add51;
output 	Add41;
output 	Add52;
output 	Add42;
output 	Add53;
output 	Add43;
output 	Add54;
output 	Add44;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	saved_grant_0;
output 	awready;
output 	wready;
output 	sop_enable1;
output 	burst_bytecount_6;
output 	write_cp_data_69;
output 	Add2;
output 	burst_bytecount_5;
output 	write_cp_data_68;
output 	burst_bytecount_3;
output 	write_cp_data_66;
output 	burst_bytecount_2;
output 	write_cp_data_65;
output 	burst_bytecount_4;
output 	write_cp_data_67;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_data_2;
output 	Add3;
output 	log2ceil;
output 	log2ceil1;
output 	Add1;
output 	Selector17;
input 	src_payload;
output 	out_data_4;
input 	src_payload1;
output 	out_data_3;
output 	out_data_1;
output 	Add31;
input 	src_payload2;
output 	out_data_0;
input 	src_payload3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add5~2 ;
wire \Add4~2 ;
wire \Add5~10 ;
wire \Add4~10 ;
wire \Add5~14 ;
wire \Add4~14 ;
wire \Add5~18 ;
wire \Add4~18 ;
wire \Decoder1~0_combout ;
wire \Decoder0~0_combout ;
wire \Decoder1~1_combout ;
wire \Decoder0~1_combout ;
wire \Decoder1~2_combout ;
wire \Decoder0~2_combout ;
wire \Decoder1~3_combout ;
wire \Decoder0~3_combout ;
wire \Decoder1~4_combout ;
wire \Decoder0~4_combout ;
wire \sop_enable~0_combout ;
wire \Add7~0_combout ;
wire \Add6~0_combout ;
wire \Add7~1_combout ;
wire \Add7~2_combout ;
wire \Add7~3_combout ;


Computer_System_altera_merlin_address_alignment_5 align_address_to_size(
	.h2f_lw_AWADDR_0(h2f_lw_AWADDR_0),
	.h2f_lw_AWADDR_1(h2f_lw_AWADDR_1),
	.h2f_lw_AWADDR_2(h2f_lw_AWADDR_2),
	.h2f_lw_AWADDR_3(h2f_lw_AWADDR_3),
	.h2f_lw_AWADDR_4(h2f_lw_AWADDR_4),
	.h2f_lw_AWBURST_0(h2f_lw_AWBURST_0),
	.h2f_lw_AWBURST_1(h2f_lw_AWBURST_1),
	.h2f_lw_AWLEN_3(h2f_lw_AWLEN_3),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.clk(outclk_wire_0),
	.wready(wready),
	.sop_enable(sop_enable1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.out_data_2(out_data_2),
	.log2ceil(log2ceil1),
	.Add1(Add1),
	.Selector17(Selector17),
	.src_payload(src_payload),
	.out_data_4(out_data_4),
	.src_payload1(src_payload1),
	.out_data_3(out_data_3),
	.Decoder0(\Decoder0~0_combout ),
	.Decoder01(\Decoder0~1_combout ),
	.Decoder02(\Decoder0~2_combout ),
	.Decoder03(\Decoder0~3_combout ),
	.out_data_1(out_data_1),
	.src_payload2(src_payload2),
	.Decoder04(\Decoder0~4_combout ),
	.out_data_0(out_data_0),
	.src_payload3(src_payload3));

cyclonev_lcell_comb \Add5~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add5),
	.cout(\Add5~2 ),
	.shareout());
defparam \Add5~1 .extended_lut = "off";
defparam \Add5~1 .lut_mask = 64'h00000000000000FF;
defparam \Add5~1 .shared_arith = "off";

cyclonev_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add4),
	.cout(\Add4~2 ),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h00000000000000FF;
defparam \Add4~1 .shared_arith = "off";

cyclonev_lcell_comb \Add5~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add51),
	.cout(),
	.shareout());
defparam \Add5~5 .extended_lut = "off";
defparam \Add5~5 .lut_mask = 64'h00000000000000FF;
defparam \Add5~5 .shared_arith = "off";

cyclonev_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add41),
	.cout(),
	.shareout());
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h00000000000000FF;
defparam \Add4~5 .shared_arith = "off";

cyclonev_lcell_comb \Add5~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add52),
	.cout(\Add5~10 ),
	.shareout());
defparam \Add5~9 .extended_lut = "off";
defparam \Add5~9 .lut_mask = 64'h00000000000000FF;
defparam \Add5~9 .shared_arith = "off";

cyclonev_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add42),
	.cout(\Add4~10 ),
	.shareout());
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h00000000000000FF;
defparam \Add4~9 .shared_arith = "off";

cyclonev_lcell_comb \Add5~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add53),
	.cout(\Add5~14 ),
	.shareout());
defparam \Add5~13 .extended_lut = "off";
defparam \Add5~13 .lut_mask = 64'h00000000000000FF;
defparam \Add5~13 .shared_arith = "off";

cyclonev_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add43),
	.cout(\Add4~14 ),
	.shareout());
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h00000000000000FF;
defparam \Add4~13 .shared_arith = "off";

cyclonev_lcell_comb \Add5~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add54),
	.cout(\Add5~18 ),
	.shareout());
defparam \Add5~17 .extended_lut = "off";
defparam \Add5~17 .lut_mask = 64'h00000000000000FF;
defparam \Add5~17 .shared_arith = "off";

cyclonev_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder0~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add44),
	.cout(\Add4~18 ),
	.shareout());
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h00000000000000FF;
defparam \Add4~17 .shared_arith = "off";

cyclonev_lcell_comb \awready~0 (
	.dataa(!h2f_lw_AWVALID_0),
	.datab(!h2f_lw_WLAST_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(!nxt_in_ready),
	.datae(!nxt_in_ready1),
	.dataf(!saved_grant_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(awready),
	.sumout(),
	.cout(),
	.shareout());
defparam \awready~0 .extended_lut = "off";
defparam \awready~0 .lut_mask = 64'h0000000000010101;
defparam \awready~0 .shared_arith = "off";

cyclonev_lcell_comb \wready~0 (
	.dataa(!h2f_lw_AWVALID_0),
	.datab(!h2f_lw_WVALID_0),
	.datac(!nxt_in_ready),
	.datad(!nxt_in_ready1),
	.datae(!saved_grant_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(wready),
	.sumout(),
	.cout(),
	.shareout());
defparam \wready~0 .extended_lut = "off";
defparam \wready~0 .lut_mask = 64'h0000011100000111;
defparam \wready~0 .shared_arith = "off";

dffeas sop_enable(
	.clk(outclk_wire_0),
	.d(\sop_enable~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(sop_enable1),
	.prn(vcc));
defparam sop_enable.is_wysiwyg = "true";
defparam sop_enable.power_up = "low";

dffeas \burst_bytecount[6] (
	.clk(outclk_wire_0),
	.d(\Add7~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_6),
	.prn(vcc));
defparam \burst_bytecount[6] .is_wysiwyg = "true";
defparam \burst_bytecount[6] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[69]~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!sop_enable1),
	.datac(!burst_bytecount_6),
	.datad(!\Add6~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_69),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[69]~0 .extended_lut = "off";
defparam \write_cp_data[69]~0 .lut_mask = 64'h0347034703470347;
defparam \write_cp_data[69]~0 .shared_arith = "off";

cyclonev_lcell_comb \Add2~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~0 .extended_lut = "off";
defparam \Add2~0 .lut_mask = 64'h0101010101010101;
defparam \Add2~0 .shared_arith = "off";

dffeas \burst_bytecount[5] (
	.clk(outclk_wire_0),
	.d(\Add7~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_5),
	.prn(vcc));
defparam \burst_bytecount[5] .is_wysiwyg = "true";
defparam \burst_bytecount[5] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[68]~1 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!sop_enable1),
	.datac(!\Add6~0_combout ),
	.datad(!burst_bytecount_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_68),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[68]~1 .extended_lut = "off";
defparam \write_cp_data[68]~1 .lut_mask = 64'h487B487B487B487B;
defparam \write_cp_data[68]~1 .shared_arith = "off";

dffeas \burst_bytecount[3] (
	.clk(outclk_wire_0),
	.d(\Add7~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_3),
	.prn(vcc));
defparam \burst_bytecount[3] .is_wysiwyg = "true";
defparam \burst_bytecount[3] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[66]~2 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!sop_enable1),
	.datad(!burst_bytecount_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_66),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[66]~2 .extended_lut = "off";
defparam \write_cp_data[66]~2 .lut_mask = 64'h606F606F606F606F;
defparam \write_cp_data[66]~2 .shared_arith = "off";

dffeas \burst_bytecount[2] (
	.clk(outclk_wire_0),
	.d(write_cp_data_65),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_2),
	.prn(vcc));
defparam \burst_bytecount[2] .is_wysiwyg = "true";
defparam \burst_bytecount[2] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[65]~3 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!sop_enable1),
	.datac(!burst_bytecount_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_65),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[65]~3 .extended_lut = "off";
defparam \write_cp_data[65]~3 .lut_mask = 64'h7474747474747474;
defparam \write_cp_data[65]~3 .shared_arith = "off";

dffeas \burst_bytecount[4] (
	.clk(outclk_wire_0),
	.d(\Add7~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(burst_bytecount_4),
	.prn(vcc));
defparam \burst_bytecount[4] .is_wysiwyg = "true";
defparam \burst_bytecount[4] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[67]~4 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!sop_enable1),
	.datae(!burst_bytecount_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_67),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[67]~4 .extended_lut = "off";
defparam \write_cp_data[67]~4 .lut_mask = 64'h1E001EFF1E001EFF;
defparam \write_cp_data[67]~4 .shared_arith = "off";

cyclonev_lcell_comb \Add3~0 (
	.dataa(!h2f_lw_ARLEN_1),
	.datab(!h2f_lw_ARLEN_2),
	.datac(!h2f_lw_ARLEN_3),
	.datad(!h2f_lw_ARSIZE_1),
	.datae(!h2f_lw_ARLEN_0),
	.dataf(!h2f_lw_ARSIZE_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~0 .extended_lut = "off";
defparam \Add3~0 .lut_mask = 64'h00700070307030F0;
defparam \Add3~0 .shared_arith = "off";

cyclonev_lcell_comb \log2ceil~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(log2ceil),
	.sumout(),
	.cout(),
	.shareout());
defparam \log2ceil~0 .extended_lut = "off";
defparam \log2ceil~0 .lut_mask = 64'h4F004F004F004F00;
defparam \log2ceil~0 .shared_arith = "off";

cyclonev_lcell_comb \log2ceil~1 (
	.dataa(!h2f_lw_AWLEN_1),
	.datab(!h2f_lw_AWLEN_2),
	.datac(!h2f_lw_AWLEN_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(log2ceil1),
	.sumout(),
	.cout(),
	.shareout());
defparam \log2ceil~1 .extended_lut = "off";
defparam \log2ceil~1 .lut_mask = 64'h7070707070707070;
defparam \log2ceil~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(!h2f_lw_AWSIZE_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h00004F0000004F00;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \Add3~1 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(!h2f_lw_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add31),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h3F007000C0FF8FFF;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~0 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~0 .extended_lut = "off";
defparam \Decoder1~0 .lut_mask = 64'h2020202020202020;
defparam \Decoder1~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'h2020202020202020;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~1 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~1 .extended_lut = "off";
defparam \Decoder1~1 .lut_mask = 64'h0808080808080808;
defparam \Decoder1~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'h0808080808080808;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~2 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~2 .extended_lut = "off";
defparam \Decoder1~2 .lut_mask = 64'h1010101010101010;
defparam \Decoder1~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~2 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~2 .extended_lut = "off";
defparam \Decoder0~2 .lut_mask = 64'h1010101010101010;
defparam \Decoder0~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~3 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~3 .extended_lut = "off";
defparam \Decoder1~3 .lut_mask = 64'h4040404040404040;
defparam \Decoder1~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~3 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~3 .extended_lut = "off";
defparam \Decoder0~3 .lut_mask = 64'h4040404040404040;
defparam \Decoder0~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~4 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~4 .extended_lut = "off";
defparam \Decoder1~4 .lut_mask = 64'h8080808080808080;
defparam \Decoder1~4 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~4 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~4 .extended_lut = "off";
defparam \Decoder0~4 .lut_mask = 64'h8080808080808080;
defparam \Decoder0~4 .shared_arith = "off";

cyclonev_lcell_comb \sop_enable~0 (
	.dataa(!h2f_lw_WLAST_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sop_enable~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sop_enable~0 .extended_lut = "off";
defparam \sop_enable~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sop_enable~0 .shared_arith = "off";

cyclonev_lcell_comb \Add7~0 (
	.dataa(!write_cp_data_69),
	.datab(!write_cp_data_68),
	.datac(!write_cp_data_66),
	.datad(!write_cp_data_65),
	.datae(!write_cp_data_67),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~0 .extended_lut = "off";
defparam \Add7~0 .lut_mask = 64'h5595555555955555;
defparam \Add7~0 .shared_arith = "off";

cyclonev_lcell_comb \Add6~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add6~0 .extended_lut = "off";
defparam \Add6~0 .lut_mask = 64'h0101010101010101;
defparam \Add6~0 .shared_arith = "off";

cyclonev_lcell_comb \Add7~1 (
	.dataa(!write_cp_data_68),
	.datab(!write_cp_data_66),
	.datac(!write_cp_data_65),
	.datad(!write_cp_data_67),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h5955595559555955;
defparam \Add7~1 .shared_arith = "off";

cyclonev_lcell_comb \Add7~2 (
	.dataa(!write_cp_data_66),
	.datab(!write_cp_data_65),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~2 .extended_lut = "off";
defparam \Add7~2 .lut_mask = 64'h6666666666666666;
defparam \Add7~2 .shared_arith = "off";

cyclonev_lcell_comb \Add7~3 (
	.dataa(!write_cp_data_66),
	.datab(!write_cp_data_65),
	.datac(!write_cp_data_67),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~3 .extended_lut = "off";
defparam \Add7~3 .lut_mask = 64'h2D2D2D2D2D2D2D2D;
defparam \Add7~3 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_address_alignment_5 (
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	clk,
	wready,
	sop_enable,
	reset,
	out_data_2,
	log2ceil,
	Add1,
	Selector17,
	src_payload,
	out_data_4,
	src_payload1,
	out_data_3,
	Decoder0,
	Decoder01,
	Decoder02,
	Decoder03,
	out_data_1,
	src_payload2,
	Decoder04,
	out_data_0,
	src_payload3)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	clk;
input 	wready;
input 	sop_enable;
input 	reset;
output 	out_data_2;
input 	log2ceil;
input 	Add1;
output 	Selector17;
input 	src_payload;
output 	out_data_4;
input 	src_payload1;
output 	out_data_3;
input 	Decoder0;
input 	Decoder01;
input 	Decoder02;
input 	Decoder03;
output 	out_data_1;
input 	src_payload2;
input 	Decoder04;
output 	out_data_0;
input 	src_payload3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add1~17_sumout ;
wire \Add0~17_sumout ;
wire \Selector20~0_combout ;
wire \address_burst[0]~q ;
wire \Add1~18 ;
wire \Add1~13_sumout ;
wire \aligned_address_bits[1]~combout ;
wire \Add0~18 ;
wire \Add0~13_sumout ;
wire \Selector19~0_combout ;
wire \address_burst[1]~q ;
wire \Add1~14 ;
wire \Add1~1_sumout ;
wire \Add0~14 ;
wire \Add0~1_sumout ;
wire \Selector18~0_combout ;
wire \address_burst[2]~q ;
wire \Add1~2 ;
wire \Add1~9_sumout ;
wire \Add0~2 ;
wire \Add0~9_sumout ;
wire \Selector17~1_combout ;
wire \address_burst[3]~q ;
wire \Add1~10 ;
wire \Add1~5_sumout ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \Selector16~0_combout ;
wire \address_burst[4]~q ;


cyclonev_lcell_comb \out_data[2]~0 (
	.dataa(!h2f_lw_AWADDR_2),
	.datab(!sop_enable),
	.datac(!\address_burst[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[2]~0 .extended_lut = "off";
defparam \out_data[2]~0 .lut_mask = 64'h4747474747474747;
defparam \out_data[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!Add1),
	.datae(!log2ceil),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector17),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~0 .extended_lut = "off";
defparam \Selector17~0 .lut_mask = 64'hA0808000A0808000;
defparam \Selector17~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[4]~1 (
	.dataa(!h2f_lw_AWADDR_4),
	.datab(!sop_enable),
	.datac(!\address_burst[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[4]~1 .extended_lut = "off";
defparam \out_data[4]~1 .lut_mask = 64'h4747474747474747;
defparam \out_data[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[3]~2 (
	.dataa(!h2f_lw_AWADDR_3),
	.datab(!sop_enable),
	.datac(!\address_burst[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[3]~2 .extended_lut = "off";
defparam \out_data[3]~2 .lut_mask = 64'h4747474747474747;
defparam \out_data[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \out_data[1]~3 (
	.dataa(!h2f_lw_AWADDR_1),
	.datab(!sop_enable),
	.datac(!\address_burst[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[1]~3 .extended_lut = "off";
defparam \out_data[1]~3 .lut_mask = 64'h4747474747474747;
defparam \out_data[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \out_data[0]~4 (
	.dataa(!h2f_lw_AWADDR_0),
	.datab(!sop_enable),
	.datac(!\address_burst[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[0]~4 .extended_lut = "off";
defparam \out_data[0]~4 .lut_mask = 64'h4747474747474747;
defparam \out_data[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[0]~q ),
	.datad(!Decoder04),
	.datae(gnd),
	.dataf(!h2f_lw_AWADDR_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(!sop_enable),
	.datab(!\address_burst[0]~q ),
	.datac(!h2f_lw_AWADDR_0),
	.datad(!Decoder04),
	.datae(gnd),
	.dataf(!Decoder04),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000EEE4000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Selector20~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\Add1~17_sumout ),
	.datad(!\Add0~17_sumout ),
	.datae(!out_data_0),
	.dataf(!src_payload3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~0 .extended_lut = "off";
defparam \Selector20~0 .lut_mask = 64'h02578ADF0055AAFF;
defparam \Selector20~0 .shared_arith = "off";

dffeas \address_burst[0] (
	.clk(clk),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\address_burst[0]~q ),
	.prn(vcc));
defparam \address_burst[0] .is_wysiwyg = "true";
defparam \address_burst[0] .power_up = "low";

cyclonev_lcell_comb \Add1~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[1]~q ),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!h2f_lw_AWADDR_1),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \aligned_address_bits[1] (
	.dataa(!h2f_lw_AWADDR_1),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aligned_address_bits[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aligned_address_bits[1] .extended_lut = "off";
defparam \aligned_address_bits[1] .lut_mask = 64'h4040404040404040;
defparam \aligned_address_bits[1] .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[1]~q ),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!\aligned_address_bits[1]~combout ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FA50000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Selector19~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\Add1~13_sumout ),
	.datad(!\Add0~13_sumout ),
	.datae(!out_data_1),
	.dataf(!src_payload2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector19~0 .extended_lut = "off";
defparam \Selector19~0 .lut_mask = 64'h02578ADF0055AAFF;
defparam \Selector19~0 .shared_arith = "off";

dffeas \address_burst[1] (
	.clk(clk),
	.d(\Selector19~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\address_burst[1]~q ),
	.prn(vcc));
defparam \address_burst[1] .is_wysiwyg = "true";
defparam \address_burst[1] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_2),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!\address_burst[2]~q ),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_2),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!\address_burst[2]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector18~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!out_data_2),
	.datad(!src_payload),
	.datae(!\Add1~1_sumout ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector18~0 .extended_lut = "off";
defparam \Selector18~0 .lut_mask = 64'h080A2A0A5D5F7F5F;
defparam \Selector18~0 .shared_arith = "off";

dffeas \address_burst[2] (
	.clk(clk),
	.d(\Selector18~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\address_burst[2]~q ),
	.prn(vcc));
defparam \address_burst[2] .is_wysiwyg = "true";
defparam \address_burst[2] .power_up = "low";

cyclonev_lcell_comb \Add1~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_3),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!\address_burst[3]~q ),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_3),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!\address_burst[3]~q ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~1 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!Selector17),
	.datad(!out_data_3),
	.datae(!\Add1~9_sumout ),
	.dataf(!\Add0~9_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~1 .extended_lut = "off";
defparam \Selector17~1 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector17~1 .shared_arith = "off";

dffeas \address_burst[3] (
	.clk(clk),
	.d(\Selector17~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\address_burst[3]~q ),
	.prn(vcc));
defparam \address_burst[3] .is_wysiwyg = "true";
defparam \address_burst[3] .power_up = "low";

cyclonev_lcell_comb \Add1~5 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_4),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!\address_burst[4]~q ),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_4),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!\address_burst[4]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!out_data_4),
	.datad(!src_payload1),
	.datae(!\Add1~5_sumout ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~0 .extended_lut = "off";
defparam \Selector16~0 .lut_mask = 64'h080A2A0A5D5F7F5F;
defparam \Selector16~0 .shared_arith = "off";

dffeas \address_burst[4] (
	.clk(clk),
	.d(\Selector16~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wready),
	.q(\address_burst[4]~q ),
	.prn(vcc));
defparam \address_burst[4] .is_wysiwyg = "true";
defparam \address_burst[4] .power_up = "low";

endmodule

module Computer_System_altera_merlin_burst_adapter_2 (
	h2f_lw_AWVALID_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	outclk_wire_0,
	saved_grant_1,
	stateST_COMP_TRANS,
	in_ready_hold,
	stateST_UNCOMP_WR_SUBBURST,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_0,
	in_data_reg_59,
	cp_ready,
	nxt_in_ready,
	local_write,
	write,
	nxt_in_ready1,
	saved_grant_0,
	r_sync_rst,
	WideOr1,
	src_payload_0,
	nxt_out_eop,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	cp_ready1,
	in_data_reg_60,
	src_data_78,
	src_data_79,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	sop_enable,
	burst_bytecount_6,
	write_cp_data_69,
	Add2,
	burst_bytecount_5,
	write_cp_data_68,
	burst_bytecount_3,
	write_cp_data_66,
	burst_bytecount_2,
	write_cp_data_65,
	burst_bytecount_4,
	write_cp_data_67,
	in_data_reg_88,
	in_data_reg_89,
	in_data_reg_90,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	src_data_88,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_3,
	out_data_2,
	src_data_72,
	out_data_4,
	src_data_74,
	out_data_3,
	src_data_73,
	in_data_reg_0,
	in_data_reg_2,
	in_data_reg_1,
	in_data_reg_14,
	in_data_reg_8,
	in_data_reg_13,
	in_data_reg_12,
	in_data_reg_11,
	in_data_reg_10,
	in_data_reg_9,
	in_data_reg_19,
	in_data_reg_18,
	in_data_reg_17,
	in_data_reg_16,
	in_data_reg_15,
	in_data_reg_26,
	in_data_reg_21,
	in_data_reg_20,
	in_data_reg_31,
	in_data_reg_30,
	in_data_reg_29,
	in_data_reg_28,
	in_data_reg_27,
	in_data_reg_25,
	in_data_reg_24,
	in_data_reg_23,
	in_data_reg_22,
	in_data_reg_7,
	in_data_reg_6,
	in_data_reg_5,
	in_data_reg_4,
	in_data_reg_3,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_data_77,
	out_data_1,
	src_data_71,
	out_data_0,
	src_data_70)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	outclk_wire_0;
input 	saved_grant_1;
output 	stateST_COMP_TRANS;
output 	in_ready_hold;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	out_valid_reg;
input 	mem_used_1;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
input 	WideOr0;
input 	wait_latency_counter_0;
output 	in_data_reg_59;
input 	cp_ready;
output 	nxt_in_ready;
input 	local_write;
input 	write;
output 	nxt_in_ready1;
input 	saved_grant_0;
input 	r_sync_rst;
input 	WideOr1;
input 	src_payload_0;
output 	nxt_out_eop;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
input 	cp_ready1;
output 	in_data_reg_60;
input 	src_data_78;
input 	src_data_79;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
input 	sop_enable;
input 	burst_bytecount_6;
input 	write_cp_data_69;
input 	Add2;
input 	burst_bytecount_5;
input 	write_cp_data_68;
input 	burst_bytecount_3;
input 	write_cp_data_66;
input 	burst_bytecount_2;
input 	write_cp_data_65;
input 	burst_bytecount_4;
input 	write_cp_data_67;
output 	in_data_reg_88;
output 	in_data_reg_89;
output 	in_data_reg_90;
output 	in_data_reg_91;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
input 	src_data_88;
input 	src_data_89;
input 	src_data_90;
input 	src_data_91;
input 	src_data_92;
input 	src_data_93;
input 	src_data_94;
input 	src_data_95;
input 	src_data_96;
input 	src_data_97;
input 	src_data_98;
input 	src_data_99;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_3;
input 	out_data_2;
input 	src_data_72;
input 	out_data_4;
input 	src_data_74;
input 	out_data_3;
input 	src_data_73;
output 	in_data_reg_0;
output 	in_data_reg_2;
output 	in_data_reg_1;
output 	in_data_reg_14;
output 	in_data_reg_8;
output 	in_data_reg_13;
output 	in_data_reg_12;
output 	in_data_reg_11;
output 	in_data_reg_10;
output 	in_data_reg_9;
output 	in_data_reg_19;
output 	in_data_reg_18;
output 	in_data_reg_17;
output 	in_data_reg_16;
output 	in_data_reg_15;
output 	in_data_reg_26;
output 	in_data_reg_21;
output 	in_data_reg_20;
output 	in_data_reg_31;
output 	in_data_reg_30;
output 	in_data_reg_29;
output 	in_data_reg_28;
output 	in_data_reg_27;
output 	in_data_reg_25;
output 	in_data_reg_24;
output 	in_data_reg_23;
output 	in_data_reg_22;
output 	in_data_reg_7;
output 	in_data_reg_6;
output 	in_data_reg_5;
output 	in_data_reg_4;
output 	in_data_reg_3;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_data_77;
input 	out_data_1;
input 	src_data_71;
input 	out_data_0;
input 	src_data_70;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altera_merlin_burst_adapter_13_1_2 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARADDR_4(h2f_lw_ARADDR_4),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.outclk_wire_0(outclk_wire_0),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_99,src_data_98,src_data_97,src_data_96,src_data_95,src_data_94,src_data_93,src_data_92,src_data_91,src_data_90,src_data_89,src_data_88,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_79,src_data_78,
src_data_77,gnd,gnd,src_data_74,src_data_73,src_data_72,src_data_71,src_data_70,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,src_data_32,src_payload18,
src_payload19,src_payload20,src_payload21,src_payload22,src_payload15,src_payload23,src_payload24,src_payload25,src_payload26,src_payload16,src_payload17,src_payload10,src_payload11,src_payload12,src_payload13,src_payload14,src_payload3,src_payload5,src_payload6,src_payload7,
src_payload8,src_payload9,src_payload4,src_payload27,src_payload28,src_payload29,src_payload30,src_payload31,src_payload1,src_payload2,src_payload}),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.in_ready_hold1(in_ready_hold),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.out_valid_reg1(out_valid_reg),
	.mem_used_1(mem_used_1),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.WideOr01(WideOr0),
	.wait_latency_counter_0(wait_latency_counter_0),
	.in_data_reg_59(in_data_reg_59),
	.cp_ready(cp_ready),
	.nxt_in_ready(nxt_in_ready),
	.local_write(local_write),
	.write(write),
	.nxt_in_ready1(nxt_in_ready1),
	.r_sync_rst(r_sync_rst),
	.WideOr1(WideOr1),
	.sink0_endofpacket(src_payload_0),
	.nxt_out_eop(nxt_out_eop),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.cp_ready1(cp_ready1),
	.in_data_reg_60(in_data_reg_60),
	.sop_enable(sop_enable),
	.burst_bytecount_6(burst_bytecount_6),
	.write_cp_data_69(write_cp_data_69),
	.Add2(Add2),
	.burst_bytecount_5(burst_bytecount_5),
	.write_cp_data_68(write_cp_data_68),
	.burst_bytecount_3(burst_bytecount_3),
	.write_cp_data_66(write_cp_data_66),
	.burst_bytecount_2(burst_bytecount_2),
	.write_cp_data_65(write_cp_data_65),
	.burst_bytecount_4(burst_bytecount_4),
	.write_cp_data_67(write_cp_data_67),
	.in_data_reg_88(in_data_reg_88),
	.in_data_reg_89(in_data_reg_89),
	.in_data_reg_90(in_data_reg_90),
	.in_data_reg_91(in_data_reg_91),
	.in_data_reg_92(in_data_reg_92),
	.in_data_reg_93(in_data_reg_93),
	.in_data_reg_94(in_data_reg_94),
	.in_data_reg_95(in_data_reg_95),
	.in_data_reg_96(in_data_reg_96),
	.in_data_reg_97(in_data_reg_97),
	.in_data_reg_98(in_data_reg_98),
	.in_data_reg_99(in_data_reg_99),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.int_nxt_addr_reg_dly_4(int_nxt_addr_reg_dly_4),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.out_data_2(out_data_2),
	.out_data_4(out_data_4),
	.out_data_3(out_data_3),
	.in_data_reg_0(in_data_reg_0),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_31(in_data_reg_31),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_24(in_data_reg_24),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_3(in_data_reg_3),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0));

endmodule

module Computer_System_altera_merlin_burst_adapter_13_1_2 (
	h2f_lw_AWVALID_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	outclk_wire_0,
	sink0_data,
	stateST_COMP_TRANS,
	in_ready_hold1,
	stateST_UNCOMP_WR_SUBBURST,
	out_valid_reg1,
	mem_used_1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr01,
	wait_latency_counter_0,
	in_data_reg_59,
	cp_ready,
	nxt_in_ready,
	local_write,
	write,
	nxt_in_ready1,
	r_sync_rst,
	WideOr1,
	sink0_endofpacket,
	nxt_out_eop,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	cp_ready1,
	in_data_reg_60,
	sop_enable,
	burst_bytecount_6,
	write_cp_data_69,
	Add2,
	burst_bytecount_5,
	write_cp_data_68,
	burst_bytecount_3,
	write_cp_data_66,
	burst_bytecount_2,
	write_cp_data_65,
	burst_bytecount_4,
	write_cp_data_67,
	in_data_reg_88,
	in_data_reg_89,
	in_data_reg_90,
	in_data_reg_91,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_3,
	out_data_2,
	out_data_4,
	out_data_3,
	in_data_reg_0,
	in_data_reg_2,
	in_data_reg_1,
	in_data_reg_14,
	in_data_reg_8,
	in_data_reg_13,
	in_data_reg_12,
	in_data_reg_11,
	in_data_reg_10,
	in_data_reg_9,
	in_data_reg_19,
	in_data_reg_18,
	in_data_reg_17,
	in_data_reg_16,
	in_data_reg_15,
	in_data_reg_26,
	in_data_reg_21,
	in_data_reg_20,
	in_data_reg_31,
	in_data_reg_30,
	in_data_reg_29,
	in_data_reg_28,
	in_data_reg_27,
	in_data_reg_25,
	in_data_reg_24,
	in_data_reg_23,
	in_data_reg_22,
	in_data_reg_7,
	in_data_reg_6,
	in_data_reg_5,
	in_data_reg_4,
	in_data_reg_3,
	out_data_1,
	out_data_0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	outclk_wire_0;
input 	[124:0] sink0_data;
output 	stateST_COMP_TRANS;
output 	in_ready_hold1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	out_valid_reg1;
input 	mem_used_1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
input 	WideOr01;
input 	wait_latency_counter_0;
output 	in_data_reg_59;
input 	cp_ready;
output 	nxt_in_ready;
input 	local_write;
input 	write;
output 	nxt_in_ready1;
input 	r_sync_rst;
input 	WideOr1;
input 	sink0_endofpacket;
output 	nxt_out_eop;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
input 	cp_ready1;
output 	in_data_reg_60;
input 	sop_enable;
input 	burst_bytecount_6;
input 	write_cp_data_69;
input 	Add2;
input 	burst_bytecount_5;
input 	write_cp_data_68;
input 	burst_bytecount_3;
input 	write_cp_data_66;
input 	burst_bytecount_2;
input 	write_cp_data_65;
input 	burst_bytecount_4;
input 	write_cp_data_67;
output 	in_data_reg_88;
output 	in_data_reg_89;
output 	in_data_reg_90;
output 	in_data_reg_91;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	int_nxt_addr_reg_dly_2;
output 	int_nxt_addr_reg_dly_4;
output 	int_nxt_addr_reg_dly_3;
input 	out_data_2;
input 	out_data_4;
input 	out_data_3;
output 	in_data_reg_0;
output 	in_data_reg_2;
output 	in_data_reg_1;
output 	in_data_reg_14;
output 	in_data_reg_8;
output 	in_data_reg_13;
output 	in_data_reg_12;
output 	in_data_reg_11;
output 	in_data_reg_10;
output 	in_data_reg_9;
output 	in_data_reg_19;
output 	in_data_reg_18;
output 	in_data_reg_17;
output 	in_data_reg_16;
output 	in_data_reg_15;
output 	in_data_reg_26;
output 	in_data_reg_21;
output 	in_data_reg_20;
output 	in_data_reg_31;
output 	in_data_reg_30;
output 	in_data_reg_29;
output 	in_data_reg_28;
output 	in_data_reg_27;
output 	in_data_reg_25;
output 	in_data_reg_24;
output 	in_data_reg_23;
output 	in_data_reg_22;
output 	in_data_reg_7;
output 	in_data_reg_6;
output 	in_data_reg_5;
output 	in_data_reg_4;
output 	in_data_reg_3;
input 	out_data_1;
input 	out_data_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \in_valid~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideOr0~combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \Selector3~0_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[2]~6_combout ;
wire \d0_int_bytes_remaining[2]~7_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~4_combout ;
wire \d0_int_bytes_remaining[3]~5_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~8_combout ;
wire \d0_int_bytes_remaining[4]~9_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~2_combout ;
wire \d0_int_bytes_remaining[5]~3_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[6]~0_combout ;
wire \d0_int_bytes_remaining[6]~1_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \WideNor0~0_combout ;
wire \WideNor0~1_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \LessThan0~0_combout ;
wire \in_eop_reg~q ;
wire \d0_int_nxt_addr[2]~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[1]~q ;
wire \in_size_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~17_sumout ;
wire \d0_int_nxt_addr[0]~9_combout ;
wire \d0_int_nxt_addr[0]~8_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~18 ;
wire \Add0~13_sumout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \d0_int_nxt_addr[1]~6_combout ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~14 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \d0_int_nxt_addr[4]~2_combout ;
wire \in_burstwrap_reg[4]~q ;
wire \nxt_addr[4]~combout ;
wire \int_nxt_addr_reg[4]~q ;
wire \ShiftLeft0~5_combout ;
wire \int_byte_cnt_narrow_reg[4]~0_combout ;
wire \int_byte_cnt_narrow_reg[4]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \Add0~2 ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[4]~3_combout ;
wire \d0_int_nxt_addr[3]~4_combout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[3]~5_combout ;


Computer_System_altera_merlin_address_alignment_6 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_77(sink0_data[77]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

dffeas \state.ST_COMP_TRANS (
	.clk(outclk_wire_0),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas in_ready_hold(
	.clk(outclk_wire_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_ready_hold1),
	.prn(vcc));
defparam in_ready_hold.is_wysiwyg = "true";
defparam in_ready_hold.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(outclk_wire_0),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

dffeas out_valid_reg(
	.clk(outclk_wire_0),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(outclk_wire_0),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[59] (
	.clk(outclk_wire_0),
	.d(sink0_data[59]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_59),
	.prn(vcc));
defparam \in_data_reg[59] .is_wysiwyg = "true";
defparam \in_data_reg[59] .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_ready_hold1),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!stateST_UNCOMP_WR_SUBBURST),
	.datae(!\load_next_out_cmd~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h20002AAA20002AAA;
defparam \nxt_in_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!write),
	.datad(gnd),
	.datae(!\new_burst_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h4444454544444545;
defparam \nxt_in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!write),
	.datac(!\in_eop_reg~q ),
	.datad(!\new_burst_reg~q ),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h0A1B4E5F0A1B4E5F;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(outclk_wire_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(outclk_wire_0),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[60] (
	.clk(outclk_wire_0),
	.d(sink0_data[60]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_60),
	.prn(vcc));
defparam \in_data_reg[60] .is_wysiwyg = "true";
defparam \in_data_reg[60] .power_up = "low";

dffeas \in_data_reg[88] (
	.clk(outclk_wire_0),
	.d(sink0_data[88]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_88),
	.prn(vcc));
defparam \in_data_reg[88] .is_wysiwyg = "true";
defparam \in_data_reg[88] .power_up = "low";

dffeas \in_data_reg[89] (
	.clk(outclk_wire_0),
	.d(sink0_data[89]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_89),
	.prn(vcc));
defparam \in_data_reg[89] .is_wysiwyg = "true";
defparam \in_data_reg[89] .power_up = "low";

dffeas \in_data_reg[90] (
	.clk(outclk_wire_0),
	.d(sink0_data[90]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_90),
	.prn(vcc));
defparam \in_data_reg[90] .is_wysiwyg = "true";
defparam \in_data_reg[90] .power_up = "low";

dffeas \in_data_reg[91] (
	.clk(outclk_wire_0),
	.d(sink0_data[91]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_91),
	.prn(vcc));
defparam \in_data_reg[91] .is_wysiwyg = "true";
defparam \in_data_reg[91] .power_up = "low";

dffeas \in_data_reg[92] (
	.clk(outclk_wire_0),
	.d(sink0_data[92]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_92),
	.prn(vcc));
defparam \in_data_reg[92] .is_wysiwyg = "true";
defparam \in_data_reg[92] .power_up = "low";

dffeas \in_data_reg[93] (
	.clk(outclk_wire_0),
	.d(sink0_data[93]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_93),
	.prn(vcc));
defparam \in_data_reg[93] .is_wysiwyg = "true";
defparam \in_data_reg[93] .power_up = "low";

dffeas \in_data_reg[94] (
	.clk(outclk_wire_0),
	.d(sink0_data[94]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_94),
	.prn(vcc));
defparam \in_data_reg[94] .is_wysiwyg = "true";
defparam \in_data_reg[94] .power_up = "low";

dffeas \in_data_reg[95] (
	.clk(outclk_wire_0),
	.d(sink0_data[95]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_95),
	.prn(vcc));
defparam \in_data_reg[95] .is_wysiwyg = "true";
defparam \in_data_reg[95] .power_up = "low";

dffeas \in_data_reg[96] (
	.clk(outclk_wire_0),
	.d(sink0_data[96]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_96),
	.prn(vcc));
defparam \in_data_reg[96] .is_wysiwyg = "true";
defparam \in_data_reg[96] .power_up = "low";

dffeas \in_data_reg[97] (
	.clk(outclk_wire_0),
	.d(sink0_data[97]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_97),
	.prn(vcc));
defparam \in_data_reg[97] .is_wysiwyg = "true";
defparam \in_data_reg[97] .power_up = "low";

dffeas \in_data_reg[98] (
	.clk(outclk_wire_0),
	.d(sink0_data[98]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_98),
	.prn(vcc));
defparam \in_data_reg[98] .is_wysiwyg = "true";
defparam \in_data_reg[98] .power_up = "low";

dffeas \in_data_reg[99] (
	.clk(outclk_wire_0),
	.d(sink0_data[99]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_99),
	.prn(vcc));
defparam \in_data_reg[99] .is_wysiwyg = "true";
defparam \in_data_reg[99] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[4] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[4]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_4),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[4] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[4] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \in_data_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \in_data_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_2),
	.prn(vcc));
defparam \in_data_reg[2] .is_wysiwyg = "true";
defparam \in_data_reg[2] .power_up = "low";

dffeas \in_data_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_1),
	.prn(vcc));
defparam \in_data_reg[1] .is_wysiwyg = "true";
defparam \in_data_reg[1] .power_up = "low";

dffeas \in_data_reg[14] (
	.clk(outclk_wire_0),
	.d(sink0_data[14]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_14),
	.prn(vcc));
defparam \in_data_reg[14] .is_wysiwyg = "true";
defparam \in_data_reg[14] .power_up = "low";

dffeas \in_data_reg[8] (
	.clk(outclk_wire_0),
	.d(sink0_data[8]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_8),
	.prn(vcc));
defparam \in_data_reg[8] .is_wysiwyg = "true";
defparam \in_data_reg[8] .power_up = "low";

dffeas \in_data_reg[13] (
	.clk(outclk_wire_0),
	.d(sink0_data[13]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_13),
	.prn(vcc));
defparam \in_data_reg[13] .is_wysiwyg = "true";
defparam \in_data_reg[13] .power_up = "low";

dffeas \in_data_reg[12] (
	.clk(outclk_wire_0),
	.d(sink0_data[12]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_12),
	.prn(vcc));
defparam \in_data_reg[12] .is_wysiwyg = "true";
defparam \in_data_reg[12] .power_up = "low";

dffeas \in_data_reg[11] (
	.clk(outclk_wire_0),
	.d(sink0_data[11]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_11),
	.prn(vcc));
defparam \in_data_reg[11] .is_wysiwyg = "true";
defparam \in_data_reg[11] .power_up = "low";

dffeas \in_data_reg[10] (
	.clk(outclk_wire_0),
	.d(sink0_data[10]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_10),
	.prn(vcc));
defparam \in_data_reg[10] .is_wysiwyg = "true";
defparam \in_data_reg[10] .power_up = "low";

dffeas \in_data_reg[9] (
	.clk(outclk_wire_0),
	.d(sink0_data[9]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_9),
	.prn(vcc));
defparam \in_data_reg[9] .is_wysiwyg = "true";
defparam \in_data_reg[9] .power_up = "low";

dffeas \in_data_reg[19] (
	.clk(outclk_wire_0),
	.d(sink0_data[19]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_19),
	.prn(vcc));
defparam \in_data_reg[19] .is_wysiwyg = "true";
defparam \in_data_reg[19] .power_up = "low";

dffeas \in_data_reg[18] (
	.clk(outclk_wire_0),
	.d(sink0_data[18]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_18),
	.prn(vcc));
defparam \in_data_reg[18] .is_wysiwyg = "true";
defparam \in_data_reg[18] .power_up = "low";

dffeas \in_data_reg[17] (
	.clk(outclk_wire_0),
	.d(sink0_data[17]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_17),
	.prn(vcc));
defparam \in_data_reg[17] .is_wysiwyg = "true";
defparam \in_data_reg[17] .power_up = "low";

dffeas \in_data_reg[16] (
	.clk(outclk_wire_0),
	.d(sink0_data[16]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_16),
	.prn(vcc));
defparam \in_data_reg[16] .is_wysiwyg = "true";
defparam \in_data_reg[16] .power_up = "low";

dffeas \in_data_reg[15] (
	.clk(outclk_wire_0),
	.d(sink0_data[15]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_15),
	.prn(vcc));
defparam \in_data_reg[15] .is_wysiwyg = "true";
defparam \in_data_reg[15] .power_up = "low";

dffeas \in_data_reg[26] (
	.clk(outclk_wire_0),
	.d(sink0_data[26]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_26),
	.prn(vcc));
defparam \in_data_reg[26] .is_wysiwyg = "true";
defparam \in_data_reg[26] .power_up = "low";

dffeas \in_data_reg[21] (
	.clk(outclk_wire_0),
	.d(sink0_data[21]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_21),
	.prn(vcc));
defparam \in_data_reg[21] .is_wysiwyg = "true";
defparam \in_data_reg[21] .power_up = "low";

dffeas \in_data_reg[20] (
	.clk(outclk_wire_0),
	.d(sink0_data[20]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_20),
	.prn(vcc));
defparam \in_data_reg[20] .is_wysiwyg = "true";
defparam \in_data_reg[20] .power_up = "low";

dffeas \in_data_reg[31] (
	.clk(outclk_wire_0),
	.d(sink0_data[31]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_31),
	.prn(vcc));
defparam \in_data_reg[31] .is_wysiwyg = "true";
defparam \in_data_reg[31] .power_up = "low";

dffeas \in_data_reg[30] (
	.clk(outclk_wire_0),
	.d(sink0_data[30]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_30),
	.prn(vcc));
defparam \in_data_reg[30] .is_wysiwyg = "true";
defparam \in_data_reg[30] .power_up = "low";

dffeas \in_data_reg[29] (
	.clk(outclk_wire_0),
	.d(sink0_data[29]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_29),
	.prn(vcc));
defparam \in_data_reg[29] .is_wysiwyg = "true";
defparam \in_data_reg[29] .power_up = "low";

dffeas \in_data_reg[28] (
	.clk(outclk_wire_0),
	.d(sink0_data[28]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_28),
	.prn(vcc));
defparam \in_data_reg[28] .is_wysiwyg = "true";
defparam \in_data_reg[28] .power_up = "low";

dffeas \in_data_reg[27] (
	.clk(outclk_wire_0),
	.d(sink0_data[27]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_27),
	.prn(vcc));
defparam \in_data_reg[27] .is_wysiwyg = "true";
defparam \in_data_reg[27] .power_up = "low";

dffeas \in_data_reg[25] (
	.clk(outclk_wire_0),
	.d(sink0_data[25]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_25),
	.prn(vcc));
defparam \in_data_reg[25] .is_wysiwyg = "true";
defparam \in_data_reg[25] .power_up = "low";

dffeas \in_data_reg[24] (
	.clk(outclk_wire_0),
	.d(sink0_data[24]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_24),
	.prn(vcc));
defparam \in_data_reg[24] .is_wysiwyg = "true";
defparam \in_data_reg[24] .power_up = "low";

dffeas \in_data_reg[23] (
	.clk(outclk_wire_0),
	.d(sink0_data[23]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_23),
	.prn(vcc));
defparam \in_data_reg[23] .is_wysiwyg = "true";
defparam \in_data_reg[23] .power_up = "low";

dffeas \in_data_reg[22] (
	.clk(outclk_wire_0),
	.d(sink0_data[22]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_22),
	.prn(vcc));
defparam \in_data_reg[22] .is_wysiwyg = "true";
defparam \in_data_reg[22] .power_up = "low";

dffeas \in_data_reg[7] (
	.clk(outclk_wire_0),
	.d(sink0_data[7]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_7),
	.prn(vcc));
defparam \in_data_reg[7] .is_wysiwyg = "true";
defparam \in_data_reg[7] .power_up = "low";

dffeas \in_data_reg[6] (
	.clk(outclk_wire_0),
	.d(sink0_data[6]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_6),
	.prn(vcc));
defparam \in_data_reg[6] .is_wysiwyg = "true";
defparam \in_data_reg[6] .power_up = "low";

dffeas \in_data_reg[5] (
	.clk(outclk_wire_0),
	.d(sink0_data[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_5),
	.prn(vcc));
defparam \in_data_reg[5] .is_wysiwyg = "true";
defparam \in_data_reg[5] .power_up = "low";

dffeas \in_data_reg[4] (
	.clk(outclk_wire_0),
	.d(sink0_data[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_4),
	.prn(vcc));
defparam \in_data_reg[4] .is_wysiwyg = "true";
defparam \in_data_reg[4] .power_up = "low";

dffeas \in_data_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_3),
	.prn(vcc));
defparam \in_data_reg[3] .is_wysiwyg = "true";
defparam \in_data_reg[3] .power_up = "low";

cyclonev_lcell_comb in_valid(
	.dataa(!in_ready_hold1),
	.datab(!WideOr1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h1111111111111111;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[60]),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[59]),
	.datad(!\in_valid~combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h005FCCFF005FCCFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!mem_used_1),
	.datac(!WideOr01),
	.datad(!wait_latency_counter_0),
	.datae(!in_data_reg_59),
	.dataf(!cp_ready),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hEAEAEAEAEAEEEEEA;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(outclk_wire_0),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!h2f_lw_AWVALID_0),
	.datab(!h2f_lw_WVALID_0),
	.datac(!in_ready_hold1),
	.datad(!sink0_data[59]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h0001000100010001;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!nxt_out_eop),
	.datad(!\state.ST_IDLE~q ),
	.datae(!\Selector2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0000FF070000FF07;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!mem_used_1),
	.datac(!WideOr01),
	.datad(!wait_latency_counter_0),
	.datae(!local_write),
	.dataf(!cp_ready),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h4040404040444440;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_uncomp_byte_cnt_reg_5),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!\Add4~0_combout ),
	.datae(!out_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .lut_mask = 64'h379D3298379D3298;
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_uncomp_byte_cnt_reg_4),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(!out_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .lut_mask = 64'h33D7337733823322;
defparam \nxt_uncomp_subburst_byte_cnt[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!out_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .lut_mask = 64'h3D3738323D373832;
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_uncomp_byte_cnt_reg_5),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!\Add4~0_combout ),
	.datae(!out_byte_cnt_reg_2),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .lut_mask = 64'h058D0088FF77FA72;
defparam \nxt_uncomp_subburst_byte_cnt[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h3D2C3D2C3D2C3D2C;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[4]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[6]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!\Selector2~1_combout ),
	.datab(!sink0_data[60]),
	.datac(!\in_valid~combout ),
	.datad(!\WideOr0~combout ),
	.datae(!nxt_out_eop),
	.dataf(!\state.ST_UNCOMP_TRANS~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "on";
defparam \Selector2~2 .lut_mask = 64'h4F444444FF444C4C;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(outclk_wire_0),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!nxt_out_eop),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h0000AA800000AA80;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!sink0_data[60]),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[59]),
	.datae(!\in_valid~combout ),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3030777530303330;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!nxt_out_eop),
	.datad(!\WideOr0~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h0070007000700070;
defparam \Selector3~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[6]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~6 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!write_cp_data_65),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~6 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~7 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~7 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~7 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[2]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~4 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!write_cp_data_66),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~4 .lut_mask = 64'h060606FF060606FF;
defparam \d0_int_bytes_remaining[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~5 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(!\d0_int_bytes_remaining[3]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~5 .lut_mask = 64'h280A7D5F280A7D5F;
defparam \d0_int_bytes_remaining[3]~5 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[4]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h9CCC9CCC9CCC9CCC;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~8 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!sink0_data[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~8 .lut_mask = 64'h001E001E001E001E;
defparam \d0_int_bytes_remaining[4]~8 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~9 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[59]),
	.datac(!\Add1~1_combout ),
	.datad(!write_cp_data_67),
	.datae(!\d0_int_bytes_remaining[4]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~9 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~9 .lut_mask = 64'hA0B1F5F5A0B1F5F5;
defparam \d0_int_bytes_remaining[4]~9 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[4]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[4]~q ),
	.datac(!\int_bytes_remaining_reg[3]~q ),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h4000400040004000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~2 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!Add2),
	.datae(!write_cp_data_68),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~2 .lut_mask = 64'h11221F2F11221F2F;
defparam \d0_int_bytes_remaining[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~3 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(outclk_wire_0),
	.d(\d0_int_bytes_remaining[5]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~0 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!write_cp_data_69),
	.datae(!Add2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~0 .lut_mask = 64'h000F111F000F111F;
defparam \d0_int_bytes_remaining[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[6]~q ),
	.datac(!\int_bytes_remaining_reg[5]~q ),
	.datad(!\Add1~0_combout ),
	.datae(!\d0_int_bytes_remaining[6]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~1 .lut_mask = 64'h228277D7228277D7;
defparam \d0_int_bytes_remaining[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[6]~1_combout ),
	.datac(!\d0_int_bytes_remaining[5]~3_combout ),
	.datad(!\d0_int_bytes_remaining[3]~5_combout ),
	.datae(!\d0_int_bytes_remaining[2]~7_combout ),
	.dataf(!\d0_int_bytes_remaining[4]~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAAAAEAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(outclk_wire_0),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sop_enable),
	.datab(!burst_bytecount_6),
	.datac(!burst_bytecount_5),
	.datad(!burst_bytecount_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h4000400040004000;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \WideNor0~1 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!burst_bytecount_3),
	.datad(!burst_bytecount_2),
	.datae(!\WideNor0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~1 .extended_lut = "off";
defparam \WideNor0~1 .lut_mask = 64'h8888A8888888A888;
defparam \WideNor0~1 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!nxt_in_ready),
	.datab(!nxt_in_ready1),
	.datac(!\in_valid~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0707070707070707;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(outclk_wire_0),
	.d(\WideNor0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!mem_used_1),
	.datac(!\new_burst_reg~q ),
	.datad(!\in_bytecount_reg_zero~q ),
	.datae(!\in_valid~combout ),
	.dataf(!cp_ready1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h5500FFFF5140FFFF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[78]),
	.datab(!sink0_data[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(outclk_wire_0),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~0 (
	.dataa(!h2f_lw_ARADDR_2),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~0 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[2]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[72]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[72]),
	.datac(!\in_burstwrap_reg[2]~q ),
	.datad(!\d0_int_nxt_addr[2]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

dffeas \in_size_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[77]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[78]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(outclk_wire_0),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[79]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h10BA101010BA1010;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[79]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \in_burstwrap_reg[0] (
	.clk(outclk_wire_0),
	.d(sink0_data[70]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[70]),
	.datac(!\in_burstwrap_reg[0]~q ),
	.datad(!\d0_int_nxt_addr[0]~8_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(outclk_wire_0),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~9 (
	.dataa(!h2f_lw_ARADDR_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~9 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~9 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~9 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~8 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\align_address_to_size|LessThan0~0_combout ),
	.datac(!\int_nxt_addr_reg[0]~q ),
	.datad(!\Add0~17_sumout ),
	.datae(!\in_burstwrap_reg[0]~q ),
	.dataf(!\d0_int_nxt_addr[0]~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~8 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~8 .lut_mask = 64'h0A0A0AAA1B1B1BBB;
defparam \d0_int_nxt_addr[0]~8 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[0]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(outclk_wire_0),
	.d(sink0_data[71]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[71]),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~6 (
	.dataa(!h2f_lw_ARADDR_1),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~6 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~6 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\int_nxt_addr_reg[1]~q ),
	.datad(!\in_burstwrap_reg[1]~q ),
	.datae(!\d0_int_nxt_addr[1]~6_combout ),
	.dataf(!\ShiftLeft0~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h0A2A0A2A0A2A5F7F;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(outclk_wire_0),
	.d(\d0_int_nxt_addr[1]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\d0_int_nxt_addr[2]~0_combout ),
	.datac(!\int_nxt_addr_reg[2]~q ),
	.datad(!\Add0~1_sumout ),
	.datae(gnd),
	.dataf(!\in_burstwrap_reg[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'h1B1B1B1B1BBB1BBB;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[4]~2 (
	.dataa(!h2f_lw_ARADDR_4),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[4]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[4]~2 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[4]~2 .shared_arith = "off";

dffeas \in_burstwrap_reg[4] (
	.clk(outclk_wire_0),
	.d(sink0_data[74]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[4]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[4] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[4] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[4] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[74]),
	.datac(!\in_burstwrap_reg[4]~q ),
	.datad(!\d0_int_nxt_addr[4]~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[4] .extended_lut = "off";
defparam \nxt_addr[4] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[4] .shared_arith = "off";

dffeas \int_nxt_addr_reg[4] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[4]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[4]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[4] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[4] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~5 (
	.dataa(!\in_size_reg[0]~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[77]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\new_burst_reg~q ),
	.dataf(!sink0_data[79]),
	.datag(!\in_size_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~5 .extended_lut = "on";
defparam \ShiftLeft0~5 .lut_mask = 64'hFF5FFFFFFF5F3F3F;
defparam \ShiftLeft0~5 .shared_arith = "off";

cyclonev_lcell_comb \int_byte_cnt_narrow_reg[4]~0 (
	.dataa(!\ShiftLeft0~5_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_byte_cnt_narrow_reg[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_byte_cnt_narrow_reg[4]~0 .extended_lut = "off";
defparam \int_byte_cnt_narrow_reg[4]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \int_byte_cnt_narrow_reg[4]~0 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[4] (
	.clk(outclk_wire_0),
	.d(\int_byte_cnt_narrow_reg[4]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[4]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[4] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[4] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(outclk_wire_0),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_4),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[4]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[4]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\d0_int_nxt_addr[4]~2_combout ),
	.datac(!\int_nxt_addr_reg[4]~q ),
	.datad(!\Add0~5_sumout ),
	.datae(gnd),
	.dataf(!\in_burstwrap_reg[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[4]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[4]~3 .lut_mask = 64'h1B1B1B1B1BBB1BBB;
defparam \d0_int_nxt_addr[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~4 (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~4 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[3]~4 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(outclk_wire_0),
	.d(sink0_data[73]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[73]),
	.datac(!\in_burstwrap_reg[3]~q ),
	.datad(!\d0_int_nxt_addr[3]~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(outclk_wire_0),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~5 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\d0_int_nxt_addr[3]~4_combout ),
	.datac(!\int_nxt_addr_reg[3]~q ),
	.datad(!\Add0~9_sumout ),
	.datae(gnd),
	.dataf(!\in_burstwrap_reg[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~5 .lut_mask = 64'h1B1B1B1B1BBB1BBB;
defparam \d0_int_nxt_addr[3]~5 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_address_alignment_6 (
	new_burst_reg,
	src_data_77,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_77;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_77),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_slave_agent_2 (
	outclk_wire_0,
	stateST_COMP_TRANS,
	in_ready_hold,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_0,
	in_data_reg_59,
	wait_latency_counter_1,
	cp_ready,
	local_write1,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_112_0,
	mem_used_01,
	always0,
	mem_57_0,
	mem_113_0,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat,
	source_endofpacket,
	r_sync_rst,
	cp_ready1,
	WideOr01,
	in_data_reg_60,
	m0_write1,
	m0_read)/* synthesis synthesis_greybox=0 */;
input 	outclk_wire_0;
input 	stateST_COMP_TRANS;
input 	in_ready_hold;
input 	out_valid_reg;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_0;
input 	in_data_reg_59;
input 	wait_latency_counter_1;
output 	cp_ready;
output 	local_write1;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_112_0;
input 	mem_used_01;
output 	always0;
input 	mem_57_0;
input 	mem_113_0;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat;
output 	source_endofpacket;
input 	r_sync_rst;
output 	cp_ready1;
input 	WideOr01;
input 	in_data_reg_60;
output 	m0_write1;
output 	m0_read;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cp_ready~1_combout ;


Computer_System_altera_merlin_burst_uncompressor_4 uncompressor(
	.clk(outclk_wire_0),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.mem_used_0(mem_used_0),
	.mem_112_0(mem_112_0),
	.mem_used_01(mem_used_01),
	.always0(always0),
	.mem_57_0(mem_57_0),
	.mem_113_0(mem_113_0),
	.mem_69_0(mem_69_0),
	.mem_68_0(mem_68_0),
	.mem_67_0(mem_67_0),
	.mem_66_0(mem_66_0),
	.mem_65_0(mem_65_0),
	.last_packet_beat(last_packet_beat),
	.source_endofpacket1(source_endofpacket),
	.reset(r_sync_rst),
	.WideOr0(WideOr01));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!in_ready_hold),
	.datab(!wait_latency_counter_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'h4444444444444444;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!out_valid_reg),
	.datab(!in_data_reg_59),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(local_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!in_narrow_reg),
	.datab(!\cp_ready~1_combout ),
	.datac(!wait_latency_counter_0),
	.datad(!local_write1),
	.datae(!cp_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h22222FF222222FF2;
defparam \cp_ready~2 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!local_write1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \m0_read~0 (
	.dataa(!out_valid_reg),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!in_data_reg_60),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_read),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_read~0 .extended_lut = "off";
defparam \m0_read~0 .lut_mask = 64'h0004000400040004;
defparam \m0_read~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~1 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_burst_uncompressor_4 (
	clk,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_112_0,
	mem_used_01,
	always0,
	mem_57_0,
	mem_113_0,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat,
	source_endofpacket1,
	reset,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_112_0;
input 	mem_used_01;
output 	always0;
input 	mem_57_0;
input 	mem_113_0;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat;
output 	source_endofpacket1;
input 	reset;
input 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~1_combout ;
wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[6]~q ;
wire \last_packet_beat~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \last_packet_beat~1_combout ;


cyclonev_lcell_comb \always0~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_112_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always0),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h007F007F007F007F;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!always0),
	.datab(!mem_57_0),
	.datac(!\burst_uncompress_busy~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!\last_packet_beat~0_combout ),
	.dataf(!\last_packet_beat~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3333333222222222;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb source_endofpacket(
	.dataa(!mem_113_0),
	.datab(!last_packet_beat),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_endofpacket1),
	.sumout(),
	.cout(),
	.shareout());
defparam source_endofpacket.extended_lut = "off";
defparam source_endofpacket.lut_mask = 64'h4444444444444444;
defparam source_endofpacket.shared_arith = "off";

cyclonev_lcell_comb \always0~1 (
	.dataa(!always0),
	.datab(!WideOr0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~1 .extended_lut = "off";
defparam \always0~1 .lut_mask = 64'h1111111111111111;
defparam \always0~1 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!mem_66_0),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_67_0),
	.datab(!mem_66_0),
	.datac(!mem_65_0),
	.datad(!last_packet_beat),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!last_packet_beat),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~0_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_69_0),
	.datac(!mem_68_0),
	.datad(!mem_67_0),
	.datae(!mem_66_0),
	.dataf(!mem_65_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_slave_translator_2 (
	clk,
	in_ready_hold,
	wait_latency_counter_0,
	wait_latency_counter_1,
	cp_ready,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	reset,
	m0_write,
	m0_read,
	av_readdata)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	in_ready_hold;
output 	wait_latency_counter_0;
output 	wait_latency_counter_1;
input 	cp_ready;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
input 	reset;
input 	m0_write;
input 	m0_read;
input 	[31:0] av_readdata;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \read_latency_shift_reg~0_combout ;


dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!in_ready_hold),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write),
	.datad(!wait_latency_counter_1),
	.datae(!m0_read),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h0004404400044044;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!in_ready_hold),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write),
	.datad(!wait_latency_counter_1),
	.datae(!m0_read),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0104014401040144;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!m0_write),
	.datac(!cp_ready),
	.datad(!m0_read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0006000600060006;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_mm_interconnect_1_cmd_mux (
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	outclk_wire_0,
	Add5,
	Add4,
	Add51,
	Add41,
	Add52,
	Add42,
	Add53,
	Add43,
	Add54,
	Add44,
	saved_grant_1,
	nxt_in_ready,
	nxt_in_ready1,
	sink1_ready1,
	saved_grant_0,
	r_sync_rst,
	WideOr11,
	src_payload_0,
	src_data_78,
	src_data_79,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	src_data_88,
	src_data_89,
	src_data_90,
	src_data_91,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	Add3,
	log2ceil,
	log2ceil1,
	Add1,
	Selector17,
	src_payload,
	src_data_72,
	src_payload1,
	src_data_74,
	src_data_73,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_data_77,
	Add31,
	src_payload34,
	src_data_71,
	src_payload35,
	src_data_70)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARBURST_0;
input 	h2f_lw_ARBURST_1;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWID_0;
input 	h2f_lw_AWID_1;
input 	h2f_lw_AWID_2;
input 	h2f_lw_AWID_3;
input 	h2f_lw_AWID_4;
input 	h2f_lw_AWID_5;
input 	h2f_lw_AWID_6;
input 	h2f_lw_AWID_7;
input 	h2f_lw_AWID_8;
input 	h2f_lw_AWID_9;
input 	h2f_lw_AWID_10;
input 	h2f_lw_AWID_11;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	h2f_lw_WDATA_0;
input 	h2f_lw_WDATA_1;
input 	h2f_lw_WDATA_2;
input 	h2f_lw_WDATA_3;
input 	h2f_lw_WDATA_4;
input 	h2f_lw_WDATA_5;
input 	h2f_lw_WDATA_6;
input 	h2f_lw_WDATA_7;
input 	h2f_lw_WDATA_8;
input 	h2f_lw_WDATA_9;
input 	h2f_lw_WDATA_10;
input 	h2f_lw_WDATA_11;
input 	h2f_lw_WDATA_12;
input 	h2f_lw_WDATA_13;
input 	h2f_lw_WDATA_14;
input 	h2f_lw_WDATA_15;
input 	h2f_lw_WDATA_16;
input 	h2f_lw_WDATA_17;
input 	h2f_lw_WDATA_18;
input 	h2f_lw_WDATA_19;
input 	h2f_lw_WDATA_20;
input 	h2f_lw_WDATA_21;
input 	h2f_lw_WDATA_22;
input 	h2f_lw_WDATA_23;
input 	h2f_lw_WDATA_24;
input 	h2f_lw_WDATA_25;
input 	h2f_lw_WDATA_26;
input 	h2f_lw_WDATA_27;
input 	h2f_lw_WDATA_28;
input 	h2f_lw_WDATA_29;
input 	h2f_lw_WDATA_30;
input 	h2f_lw_WDATA_31;
input 	h2f_lw_WSTRB_0;
input 	h2f_lw_WSTRB_1;
input 	h2f_lw_WSTRB_2;
input 	h2f_lw_WSTRB_3;
input 	outclk_wire_0;
input 	Add5;
input 	Add4;
input 	Add51;
input 	Add41;
input 	Add52;
input 	Add42;
input 	Add53;
input 	Add43;
input 	Add54;
input 	Add44;
output 	saved_grant_1;
input 	nxt_in_ready;
input 	nxt_in_ready1;
output 	sink1_ready1;
output 	saved_grant_0;
input 	r_sync_rst;
output 	WideOr11;
output 	src_payload_0;
output 	src_data_78;
output 	src_data_79;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
output 	src_data_88;
output 	src_data_89;
output 	src_data_90;
output 	src_data_91;
output 	src_data_92;
output 	src_data_93;
output 	src_data_94;
output 	src_data_95;
output 	src_data_96;
output 	src_data_97;
output 	src_data_98;
output 	src_data_99;
input 	Add3;
input 	log2ceil;
input 	log2ceil1;
input 	Add1;
input 	Selector17;
output 	src_payload;
output 	src_data_72;
output 	src_payload1;
output 	src_data_74;
output 	src_data_73;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
output 	src_payload33;
output 	src_data_77;
input 	Add31;
output 	src_payload34;
output 	src_data_71;
output 	src_payload35;
output 	src_data_70;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \src_data[72]~0_combout ;
wire \src_data[70]~1_combout ;
wire \src_data[72]~2_combout ;
wire \src_data[72]~3_combout ;
wire \src_data[70]~5_combout ;
wire \src_data[74]~6_combout ;
wire \src_data[74]~7_combout ;
wire \src_data[74]~8_combout ;
wire \src_data[73]~10_combout ;
wire \src_data[73]~11_combout ;
wire \src_data[71]~13_combout ;
wire \src_data[71]~14_combout ;
wire \src_data[70]~16_combout ;
wire \src_data[70]~17_combout ;


Computer_System_altera_merlin_arbitrator_4 arb(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.clk(outclk_wire_0),
	.nxt_in_ready(nxt_in_ready),
	.nxt_in_ready1(nxt_in_ready1),
	.grant_1(\arb|grant[1]~0_combout ),
	.reset(r_sync_rst),
	.WideOr1(WideOr11),
	.src_payload_0(src_payload_0),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ));

dffeas \saved_grant[1] (
	.clk(outclk_wire_0),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb sink1_ready(
	.dataa(!saved_grant_1),
	.datab(!nxt_in_ready),
	.datac(!nxt_in_ready1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink1_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam sink1_ready.extended_lut = "off";
defparam sink1_ready.lut_mask = 64'h1515151515151515;
defparam sink1_ready.shared_arith = "off";

dffeas \saved_grant[0] (
	.clk(outclk_wire_0),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb WideOr1(
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_AWVALID_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(!saved_grant_1),
	.datae(!saved_grant_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h0055035700550357;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[78] (
	.dataa(!h2f_lw_ARSIZE_1),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_78),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[78] .extended_lut = "off";
defparam \src_data[78] .lut_mask = 64'h0537053705370537;
defparam \src_data[78] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!h2f_lw_ARSIZE_2),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0537053705370537;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_lw_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_lw_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_lw_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_lw_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_data[88] (
	.dataa(!h2f_lw_ARID_0),
	.datab(!h2f_lw_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_88),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[88] .extended_lut = "off";
defparam \src_data[88] .lut_mask = 64'h0537053705370537;
defparam \src_data[88] .shared_arith = "off";

cyclonev_lcell_comb \src_data[89] (
	.dataa(!h2f_lw_ARID_1),
	.datab(!h2f_lw_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_89),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[89] .extended_lut = "off";
defparam \src_data[89] .lut_mask = 64'h0537053705370537;
defparam \src_data[89] .shared_arith = "off";

cyclonev_lcell_comb \src_data[90] (
	.dataa(!h2f_lw_ARID_2),
	.datab(!h2f_lw_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_90),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[90] .extended_lut = "off";
defparam \src_data[90] .lut_mask = 64'h0537053705370537;
defparam \src_data[90] .shared_arith = "off";

cyclonev_lcell_comb \src_data[91] (
	.dataa(!h2f_lw_ARID_3),
	.datab(!h2f_lw_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_91),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[91] .extended_lut = "off";
defparam \src_data[91] .lut_mask = 64'h0537053705370537;
defparam \src_data[91] .shared_arith = "off";

cyclonev_lcell_comb \src_data[92] (
	.dataa(!h2f_lw_ARID_4),
	.datab(!h2f_lw_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_92),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92] .extended_lut = "off";
defparam \src_data[92] .lut_mask = 64'h0537053705370537;
defparam \src_data[92] .shared_arith = "off";

cyclonev_lcell_comb \src_data[93] (
	.dataa(!h2f_lw_ARID_5),
	.datab(!h2f_lw_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_93),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[93] .extended_lut = "off";
defparam \src_data[93] .lut_mask = 64'h0537053705370537;
defparam \src_data[93] .shared_arith = "off";

cyclonev_lcell_comb \src_data[94] (
	.dataa(!h2f_lw_ARID_6),
	.datab(!h2f_lw_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_94),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94] .extended_lut = "off";
defparam \src_data[94] .lut_mask = 64'h0537053705370537;
defparam \src_data[94] .shared_arith = "off";

cyclonev_lcell_comb \src_data[95] (
	.dataa(!h2f_lw_ARID_7),
	.datab(!h2f_lw_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_95),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95] .extended_lut = "off";
defparam \src_data[95] .lut_mask = 64'h0537053705370537;
defparam \src_data[95] .shared_arith = "off";

cyclonev_lcell_comb \src_data[96] (
	.dataa(!h2f_lw_ARID_8),
	.datab(!h2f_lw_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_96),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96] .extended_lut = "off";
defparam \src_data[96] .lut_mask = 64'h0537053705370537;
defparam \src_data[96] .shared_arith = "off";

cyclonev_lcell_comb \src_data[97] (
	.dataa(!h2f_lw_ARID_9),
	.datab(!h2f_lw_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_97),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[97] .extended_lut = "off";
defparam \src_data[97] .lut_mask = 64'h0537053705370537;
defparam \src_data[97] .shared_arith = "off";

cyclonev_lcell_comb \src_data[98] (
	.dataa(!h2f_lw_ARID_10),
	.datab(!h2f_lw_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_98),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98] .extended_lut = "off";
defparam \src_data[98] .lut_mask = 64'h0537053705370537;
defparam \src_data[98] .shared_arith = "off";

cyclonev_lcell_comb \src_data[99] (
	.dataa(!h2f_lw_ARID_11),
	.datab(!h2f_lw_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_99),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99] .extended_lut = "off";
defparam \src_data[99] .lut_mask = 64'h0537053705370537;
defparam \src_data[99] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!log2ceil),
	.datad(!log2ceil1),
	.datae(!Selector17),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h0000EDB70000EDB7;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72]~4 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!\src_data[72]~2_combout ),
	.datad(!\src_data[72]~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_72),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72]~4 .extended_lut = "off";
defparam \src_data[72]~4 .lut_mask = 64'h7350735073507350;
defparam \src_data[72]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_0),
	.datac(!h2f_lw_AWSIZE_1),
	.datad(!h2f_lw_AWSIZE_2),
	.datae(!log2ceil),
	.dataf(!log2ceil1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'hEA80AA00A800A000;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~9 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!\src_data[74]~7_combout ),
	.datad(!\src_data[74]~8_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_74),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~9 .extended_lut = "off";
defparam \src_data[74]~9 .lut_mask = 64'h7350735073507350;
defparam \src_data[74]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~12 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!\src_data[73]~10_combout ),
	.datad(!\src_data[73]~11_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_73),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~12 .extended_lut = "off";
defparam \src_data[73]~12 .lut_mask = 64'h7350735073507350;
defparam \src_data[73]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_lw_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!h2f_lw_WDATA_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h1111111111111111;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!h2f_lw_WDATA_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1111111111111111;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!h2f_lw_WDATA_14),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h1111111111111111;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!h2f_lw_WDATA_8),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h1111111111111111;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!h2f_lw_WDATA_13),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h1111111111111111;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!h2f_lw_WDATA_12),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h1111111111111111;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!h2f_lw_WDATA_11),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h1111111111111111;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!h2f_lw_WDATA_10),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h1111111111111111;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!h2f_lw_WDATA_9),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h1111111111111111;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!h2f_lw_WDATA_19),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h1111111111111111;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!h2f_lw_WDATA_18),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h1111111111111111;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!h2f_lw_WDATA_17),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h1111111111111111;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!h2f_lw_WDATA_16),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h1111111111111111;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!h2f_lw_WDATA_15),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h1111111111111111;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!h2f_lw_WDATA_26),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h1111111111111111;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!h2f_lw_WDATA_21),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h1111111111111111;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!h2f_lw_WDATA_20),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h1111111111111111;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!h2f_lw_WDATA_31),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h1111111111111111;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!h2f_lw_WDATA_30),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h1111111111111111;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!h2f_lw_WDATA_29),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h1111111111111111;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!h2f_lw_WDATA_28),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h1111111111111111;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!h2f_lw_WDATA_27),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h1111111111111111;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!h2f_lw_WDATA_25),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h1111111111111111;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!h2f_lw_WDATA_24),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h1111111111111111;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!h2f_lw_WDATA_23),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h1111111111111111;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!h2f_lw_WDATA_22),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h1111111111111111;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!h2f_lw_WDATA_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h1111111111111111;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!h2f_lw_WDATA_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h1111111111111111;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!h2f_lw_WDATA_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h1111111111111111;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!h2f_lw_WDATA_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'h1111111111111111;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~33 (
	.dataa(!h2f_lw_WDATA_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~33 .extended_lut = "off";
defparam \src_payload~33 .lut_mask = 64'h1111111111111111;
defparam \src_payload~33 .shared_arith = "off";

cyclonev_lcell_comb \src_data[77] (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_77),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[77] .extended_lut = "off";
defparam \src_data[77] .lut_mask = 64'h0537053705370537;
defparam \src_data[77] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~34 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!Add1),
	.datae(!log2ceil1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~34 .extended_lut = "off";
defparam \src_payload~34 .lut_mask = 64'h8000000080000000;
defparam \src_payload~34 .shared_arith = "off";

cyclonev_lcell_comb \src_data[71]~15 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!\src_data[71]~13_combout ),
	.datad(!\src_data[71]~14_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_71),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71]~15 .extended_lut = "off";
defparam \src_data[71]~15 .lut_mask = 64'h7350735073507350;
defparam \src_data[71]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~35 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!log2ceil),
	.datac(!src_payload34),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~35 .extended_lut = "off";
defparam \src_payload~35 .lut_mask = 64'h0909090909090909;
defparam \src_payload~35 .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~18 (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!\src_data[70]~16_combout ),
	.datad(!\src_data[70]~17_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_70),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~18 .extended_lut = "off";
defparam \src_data[70]~18 .lut_mask = 64'h7350735073507350;
defparam \src_data[70]~18 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(outclk_wire_0),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready),
	.datab(!nxt_in_ready1),
	.datac(!WideOr11),
	.datad(!src_payload_0),
	.datae(!\packet_in_progress~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF0F70007F0F70007;
defparam \update_grant~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72]~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(!h2f_lw_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[72]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72]~0 .extended_lut = "off";
defparam \src_data[72]~0 .lut_mask = 64'h0F003000400080FF;
defparam \src_data[72]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~1 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_2),
	.datac(!Add3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[70]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~1 .extended_lut = "off";
defparam \src_data[70]~1 .lut_mask = 64'h8080808080808080;
defparam \src_data[70]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72]~2 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!Add5),
	.datad(!\src_data[72]~0_combout ),
	.datae(!\src_data[70]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[72]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72]~2 .extended_lut = "off";
defparam \src_data[72]~2 .lut_mask = 64'h8080A2808080A280;
defparam \src_data[72]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[72]~3 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!src_payload),
	.datad(!Add4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[72]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72]~3 .extended_lut = "off";
defparam \src_data[72]~3 .lut_mask = 64'h8A028A028A028A02;
defparam \src_data[72]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~5 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(!h2f_lw_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[70]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~5 .extended_lut = "off";
defparam \src_data[70]~5 .lut_mask = 64'h80FF0F0030004000;
defparam \src_data[70]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~6 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_2),
	.datac(!Add3),
	.datad(!\src_data[70]~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[74]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~6 .extended_lut = "off";
defparam \src_data[74]~6 .lut_mask = 64'h80E880E880E880E8;
defparam \src_data[74]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~7 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!Add51),
	.datad(!\src_data[74]~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[74]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~7 .extended_lut = "off";
defparam \src_data[74]~7 .lut_mask = 64'h80A280A280A280A2;
defparam \src_data[74]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[74]~8 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!src_payload1),
	.datad(!Add41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[74]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[74]~8 .extended_lut = "off";
defparam \src_data[74]~8 .lut_mask = 64'h8A028A028A028A02;
defparam \src_data[74]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~10 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!\src_data[70]~1_combout ),
	.datad(!Add52),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[73]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~10 .extended_lut = "off";
defparam \src_data[73]~10 .lut_mask = 64'h8A028A028A028A02;
defparam \src_data[73]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73]~11 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!Selector17),
	.datad(!Add42),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[73]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73]~11 .extended_lut = "off";
defparam \src_data[73]~11 .lut_mask = 64'h8A028A028A028A02;
defparam \src_data[73]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[71]~13 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!Add31),
	.datad(!\src_data[70]~1_combout ),
	.datae(!Add53),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[71]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71]~13 .extended_lut = "off";
defparam \src_data[71]~13 .lut_mask = 64'h88A8002088A80020;
defparam \src_data[71]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[71]~14 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!Add43),
	.datad(!src_payload34),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[71]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71]~14 .extended_lut = "off";
defparam \src_data[71]~14 .lut_mask = 64'h80A280A280A280A2;
defparam \src_data[71]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~16 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!\src_data[70]~1_combout ),
	.datad(!\src_data[70]~5_combout ),
	.datae(!Add54),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[70]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~16 .extended_lut = "off";
defparam \src_data[70]~16 .lut_mask = 64'h888A0002888A0002;
defparam \src_data[70]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[70]~17 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!Add44),
	.datad(!h2f_lw_AWSIZE_0),
	.datae(!log2ceil),
	.dataf(!src_payload34),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[70]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70]~17 .extended_lut = "off";
defparam \src_data[70]~17 .lut_mask = 64'h80808080A28080A2;
defparam \src_data[70]~17 .shared_arith = "off";

endmodule

module Computer_System_altera_merlin_arbitrator_4 (
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_WVALID_0,
	clk,
	nxt_in_ready,
	nxt_in_ready1,
	grant_1,
	reset,
	WideOr1,
	src_payload_0,
	packet_in_progress,
	grant_0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WVALID_0;
input 	clk;
input 	nxt_in_ready;
input 	nxt_in_ready1;
output 	grant_1;
input 	reset;
input 	WideOr1;
input 	src_payload_0;
input 	packet_in_progress;
output 	grant_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_AWVALID_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(!\top_priority_reg[1]~q ),
	.datae(!\top_priority_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h5455005554550055;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_AWVALID_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(!\top_priority_reg[1]~q ),
	.datae(!\top_priority_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0303000203030002;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!h2f_lw_AWVALID_0),
	.datac(!h2f_lw_WVALID_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hA8A8A8A8A8A8A8A8;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready),
	.datab(!nxt_in_ready1),
	.datac(!WideOr1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hF0F7000700000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module Computer_System_Computer_System_mm_interconnect_1_rsp_demux (
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	always0,
	mem_59_0,
	mem_57_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	always0;
input 	mem_59_0;
input 	mem_57_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src0_valid~0_combout ;


cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!always0),
	.datad(!\src0_valid~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h007F007F007F007F;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!always0),
	.datad(!\src0_valid~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F007F007F007F00;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!h2f_lw_RREADY_0),
	.datac(!\src0_valid~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3535353535353535;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!mem_59_0),
	.datab(!mem_57_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src0_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'h4444444444444444;
defparam \src0_valid~0 .shared_arith = "off";

endmodule

module Computer_System_Computer_System_Onchip_SRAM (
	q_a_0,
	q_b_0,
	q_a_1,
	q_b_1,
	q_a_2,
	q_b_2,
	q_a_3,
	q_b_3,
	q_a_4,
	q_b_4,
	q_a_5,
	q_b_5,
	q_a_6,
	q_b_6,
	q_a_7,
	q_b_7,
	q_a_8,
	q_b_8,
	q_a_9,
	q_b_9,
	q_a_10,
	q_b_10,
	q_a_11,
	q_b_11,
	q_a_12,
	q_b_12,
	q_a_13,
	q_b_13,
	q_a_14,
	q_b_14,
	q_a_15,
	q_b_15,
	q_a_16,
	q_b_16,
	q_a_17,
	q_b_17,
	q_a_18,
	q_b_18,
	q_a_19,
	q_b_19,
	q_a_20,
	q_b_20,
	q_a_21,
	q_b_21,
	q_a_22,
	q_b_22,
	q_a_23,
	q_b_23,
	q_a_24,
	q_b_24,
	q_a_25,
	q_b_25,
	q_a_26,
	q_b_26,
	q_a_27,
	q_b_27,
	q_a_28,
	q_b_28,
	q_a_29,
	q_b_29,
	q_a_30,
	q_b_30,
	q_a_31,
	q_b_31,
	outclk_wire_0,
	int_nxt_addr_reg_dly_2,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_4,
	int_nxt_addr_reg_dly_5,
	int_nxt_addr_reg_dly_6,
	int_nxt_addr_reg_dly_7,
	int_nxt_addr_reg_dly_8,
	int_nxt_addr_reg_dly_9,
	source0_data_34,
	source0_data_32,
	source0_data_33,
	source0_data_35,
	m0_write,
	r_early_rst,
	r_early_rst1,
	in_data_reg_0,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	clock_bridge_0_in_clk_clk,
	onchip_sram_s1_chipselect,
	onchip_sram_s1_write,
	onchip_sram_s1_clken,
	onchip_sram_s1_writedata_0,
	onchip_sram_s1_address_0,
	onchip_sram_s1_address_1,
	onchip_sram_s1_address_2,
	onchip_sram_s1_address_3,
	onchip_sram_s1_address_4,
	onchip_sram_s1_address_5,
	onchip_sram_s1_address_6,
	onchip_sram_s1_address_7,
	onchip_sram_s1_byteenable_0,
	onchip_sram_s1_writedata_1,
	onchip_sram_s1_writedata_2,
	onchip_sram_s1_writedata_3,
	onchip_sram_s1_writedata_4,
	onchip_sram_s1_writedata_5,
	onchip_sram_s1_writedata_6,
	onchip_sram_s1_writedata_7,
	onchip_sram_s1_writedata_8,
	onchip_sram_s1_byteenable_1,
	onchip_sram_s1_writedata_9,
	onchip_sram_s1_writedata_10,
	onchip_sram_s1_writedata_11,
	onchip_sram_s1_writedata_12,
	onchip_sram_s1_writedata_13,
	onchip_sram_s1_writedata_14,
	onchip_sram_s1_writedata_15,
	onchip_sram_s1_writedata_16,
	onchip_sram_s1_byteenable_2,
	onchip_sram_s1_writedata_17,
	onchip_sram_s1_writedata_18,
	onchip_sram_s1_writedata_19,
	onchip_sram_s1_writedata_20,
	onchip_sram_s1_writedata_21,
	onchip_sram_s1_writedata_22,
	onchip_sram_s1_writedata_23,
	onchip_sram_s1_writedata_24,
	onchip_sram_s1_byteenable_3,
	onchip_sram_s1_writedata_25,
	onchip_sram_s1_writedata_26,
	onchip_sram_s1_writedata_27,
	onchip_sram_s1_writedata_28,
	onchip_sram_s1_writedata_29,
	onchip_sram_s1_writedata_30,
	onchip_sram_s1_writedata_31)/* synthesis synthesis_greybox=0 */;
output 	q_a_0;
output 	q_b_0;
output 	q_a_1;
output 	q_b_1;
output 	q_a_2;
output 	q_b_2;
output 	q_a_3;
output 	q_b_3;
output 	q_a_4;
output 	q_b_4;
output 	q_a_5;
output 	q_b_5;
output 	q_a_6;
output 	q_b_6;
output 	q_a_7;
output 	q_b_7;
output 	q_a_8;
output 	q_b_8;
output 	q_a_9;
output 	q_b_9;
output 	q_a_10;
output 	q_b_10;
output 	q_a_11;
output 	q_b_11;
output 	q_a_12;
output 	q_b_12;
output 	q_a_13;
output 	q_b_13;
output 	q_a_14;
output 	q_b_14;
output 	q_a_15;
output 	q_b_15;
output 	q_a_16;
output 	q_b_16;
output 	q_a_17;
output 	q_b_17;
output 	q_a_18;
output 	q_b_18;
output 	q_a_19;
output 	q_b_19;
output 	q_a_20;
output 	q_b_20;
output 	q_a_21;
output 	q_b_21;
output 	q_a_22;
output 	q_b_22;
output 	q_a_23;
output 	q_b_23;
output 	q_a_24;
output 	q_b_24;
output 	q_a_25;
output 	q_b_25;
output 	q_a_26;
output 	q_b_26;
output 	q_a_27;
output 	q_b_27;
output 	q_a_28;
output 	q_b_28;
output 	q_a_29;
output 	q_b_29;
output 	q_a_30;
output 	q_b_30;
output 	q_a_31;
output 	q_b_31;
input 	outclk_wire_0;
input 	int_nxt_addr_reg_dly_2;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_4;
input 	int_nxt_addr_reg_dly_5;
input 	int_nxt_addr_reg_dly_6;
input 	int_nxt_addr_reg_dly_7;
input 	int_nxt_addr_reg_dly_8;
input 	int_nxt_addr_reg_dly_9;
input 	source0_data_34;
input 	source0_data_32;
input 	source0_data_33;
input 	source0_data_35;
input 	m0_write;
input 	r_early_rst;
input 	r_early_rst1;
input 	in_data_reg_0;
input 	in_data_reg_1;
input 	in_data_reg_2;
input 	in_data_reg_3;
input 	in_data_reg_4;
input 	in_data_reg_5;
input 	in_data_reg_6;
input 	in_data_reg_7;
input 	in_data_reg_8;
input 	in_data_reg_9;
input 	in_data_reg_10;
input 	in_data_reg_11;
input 	in_data_reg_12;
input 	in_data_reg_13;
input 	in_data_reg_14;
input 	in_data_reg_15;
input 	in_data_reg_16;
input 	in_data_reg_17;
input 	in_data_reg_18;
input 	in_data_reg_19;
input 	in_data_reg_20;
input 	in_data_reg_21;
input 	in_data_reg_22;
input 	in_data_reg_23;
input 	in_data_reg_24;
input 	in_data_reg_25;
input 	in_data_reg_26;
input 	in_data_reg_27;
input 	in_data_reg_28;
input 	in_data_reg_29;
input 	in_data_reg_30;
input 	in_data_reg_31;
input 	clock_bridge_0_in_clk_clk;
input 	onchip_sram_s1_chipselect;
input 	onchip_sram_s1_write;
input 	onchip_sram_s1_clken;
input 	onchip_sram_s1_writedata_0;
input 	onchip_sram_s1_address_0;
input 	onchip_sram_s1_address_1;
input 	onchip_sram_s1_address_2;
input 	onchip_sram_s1_address_3;
input 	onchip_sram_s1_address_4;
input 	onchip_sram_s1_address_5;
input 	onchip_sram_s1_address_6;
input 	onchip_sram_s1_address_7;
input 	onchip_sram_s1_byteenable_0;
input 	onchip_sram_s1_writedata_1;
input 	onchip_sram_s1_writedata_2;
input 	onchip_sram_s1_writedata_3;
input 	onchip_sram_s1_writedata_4;
input 	onchip_sram_s1_writedata_5;
input 	onchip_sram_s1_writedata_6;
input 	onchip_sram_s1_writedata_7;
input 	onchip_sram_s1_writedata_8;
input 	onchip_sram_s1_byteenable_1;
input 	onchip_sram_s1_writedata_9;
input 	onchip_sram_s1_writedata_10;
input 	onchip_sram_s1_writedata_11;
input 	onchip_sram_s1_writedata_12;
input 	onchip_sram_s1_writedata_13;
input 	onchip_sram_s1_writedata_14;
input 	onchip_sram_s1_writedata_15;
input 	onchip_sram_s1_writedata_16;
input 	onchip_sram_s1_byteenable_2;
input 	onchip_sram_s1_writedata_17;
input 	onchip_sram_s1_writedata_18;
input 	onchip_sram_s1_writedata_19;
input 	onchip_sram_s1_writedata_20;
input 	onchip_sram_s1_writedata_21;
input 	onchip_sram_s1_writedata_22;
input 	onchip_sram_s1_writedata_23;
input 	onchip_sram_s1_writedata_24;
input 	onchip_sram_s1_byteenable_3;
input 	onchip_sram_s1_writedata_25;
input 	onchip_sram_s1_writedata_26;
input 	onchip_sram_s1_writedata_27;
input 	onchip_sram_s1_writedata_28;
input 	onchip_sram_s1_writedata_29;
input 	onchip_sram_s1_writedata_30;
input 	onchip_sram_s1_writedata_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wren~combout ;
wire \clocken0~combout ;


Computer_System_altsyncram_1 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.clock1(outclk_wire_0),
	.address_b({int_nxt_addr_reg_dly_9,int_nxt_addr_reg_dly_8,int_nxt_addr_reg_dly_7,int_nxt_addr_reg_dly_6,int_nxt_addr_reg_dly_5,int_nxt_addr_reg_dly_4,int_nxt_addr_reg_dly_3,int_nxt_addr_reg_dly_2}),
	.byteena_b({source0_data_35,source0_data_34,source0_data_33,source0_data_32}),
	.wren_a(\wren~combout ),
	.wren_b(m0_write),
	.clocken0(\clocken0~combout ),
	.clocken1(r_early_rst1),
	.data_b({in_data_reg_31,in_data_reg_30,in_data_reg_29,in_data_reg_28,in_data_reg_27,in_data_reg_26,in_data_reg_25,in_data_reg_24,in_data_reg_23,in_data_reg_22,in_data_reg_21,in_data_reg_20,in_data_reg_19,in_data_reg_18,in_data_reg_17,in_data_reg_16,in_data_reg_15,in_data_reg_14,
in_data_reg_13,in_data_reg_12,in_data_reg_11,in_data_reg_10,in_data_reg_9,in_data_reg_8,in_data_reg_7,in_data_reg_6,in_data_reg_5,in_data_reg_4,in_data_reg_3,in_data_reg_2,in_data_reg_1,in_data_reg_0}),
	.clock0(clock_bridge_0_in_clk_clk),
	.data_a({onchip_sram_s1_writedata_31,onchip_sram_s1_writedata_30,onchip_sram_s1_writedata_29,onchip_sram_s1_writedata_28,onchip_sram_s1_writedata_27,onchip_sram_s1_writedata_26,onchip_sram_s1_writedata_25,onchip_sram_s1_writedata_24,onchip_sram_s1_writedata_23,
onchip_sram_s1_writedata_22,onchip_sram_s1_writedata_21,onchip_sram_s1_writedata_20,onchip_sram_s1_writedata_19,onchip_sram_s1_writedata_18,onchip_sram_s1_writedata_17,onchip_sram_s1_writedata_16,onchip_sram_s1_writedata_15,onchip_sram_s1_writedata_14,
onchip_sram_s1_writedata_13,onchip_sram_s1_writedata_12,onchip_sram_s1_writedata_11,onchip_sram_s1_writedata_10,onchip_sram_s1_writedata_9,onchip_sram_s1_writedata_8,onchip_sram_s1_writedata_7,onchip_sram_s1_writedata_6,onchip_sram_s1_writedata_5,
onchip_sram_s1_writedata_4,onchip_sram_s1_writedata_3,onchip_sram_s1_writedata_2,onchip_sram_s1_writedata_1,onchip_sram_s1_writedata_0}),
	.address_a({onchip_sram_s1_address_7,onchip_sram_s1_address_6,onchip_sram_s1_address_5,onchip_sram_s1_address_4,onchip_sram_s1_address_3,onchip_sram_s1_address_2,onchip_sram_s1_address_1,onchip_sram_s1_address_0}),
	.byteena_a({onchip_sram_s1_byteenable_3,onchip_sram_s1_byteenable_2,onchip_sram_s1_byteenable_1,onchip_sram_s1_byteenable_0}));

cyclonev_lcell_comb wren(
	.dataa(!onchip_sram_s1_chipselect),
	.datab(!onchip_sram_s1_write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam wren.extended_lut = "off";
defparam wren.lut_mask = 64'h1111111111111111;
defparam wren.shared_arith = "off";

cyclonev_lcell_comb clocken0(
	.dataa(!onchip_sram_s1_clken),
	.datab(!r_early_rst),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\clocken0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam clocken0.extended_lut = "off";
defparam clocken0.lut_mask = 64'h4444444444444444;
defparam clocken0.shared_arith = "off";

endmodule

module Computer_System_altsyncram_1 (
	q_a,
	q_b,
	clock1,
	address_b,
	byteena_b,
	wren_a,
	wren_b,
	clocken0,
	clocken1,
	data_b,
	clock0,
	data_a,
	address_a,
	byteena_a)/* synthesis synthesis_greybox=0 */;
output 	[31:0] q_a;
output 	[31:0] q_b;
input 	clock1;
input 	[7:0] address_b;
input 	[3:0] byteena_b;
input 	wren_a;
input 	wren_b;
input 	clocken0;
input 	clocken1;
input 	[31:0] data_b;
input 	clock0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altsyncram_1k52 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.clock1(clock1),
	.address_b({address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.byteena_b({byteena_b[3],byteena_b[2],byteena_b[1],byteena_b[0]}),
	.wren_a(wren_a),
	.wren_b(wren_b),
	.clocken0(clocken0),
	.clocken1(clocken1),
	.data_b({data_b[31],data_b[30],data_b[29],data_b[28],data_b[27],data_b[26],data_b[25],data_b[24],data_b[23],data_b[22],data_b[21],data_b[20],data_b[19],data_b[18],data_b[17],data_b[16],data_b[15],data_b[14],data_b[13],data_b[12],data_b[11],data_b[10],data_b[9],data_b[8],data_b[7],data_b[6],data_b[5],data_b[4],data_b[3],data_b[2],data_b[1],data_b[0]}),
	.clock0(clock0),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}));

endmodule

module Computer_System_altsyncram_1k52 (
	q_a,
	q_b,
	clock1,
	address_b,
	byteena_b,
	wren_a,
	wren_b,
	clocken0,
	clocken1,
	data_b,
	clock0,
	data_a,
	address_a,
	byteena_a)/* synthesis synthesis_greybox=0 */;
output 	[31:0] q_a;
output 	[31:0] q_b;
input 	clock1;
input 	[7:0] address_b;
input 	[3:0] byteena_b;
input 	wren_a;
input 	wren_b;
input 	clocken0;
input 	clocken1;
input 	[31:0] data_b;
input 	clock0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "bidir_dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 8;
defparam ram_block1a0.port_b_byte_enable_clock = "clock1";
defparam ram_block1a0.port_b_byte_enable_mask_width = 1;
defparam ram_block1a0.port_b_byte_size = 1;
defparam ram_block1a0.port_b_data_in_clock = "clock1";
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 255;
defparam ram_block1a0.port_b_logical_ram_depth = 256;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.port_b_write_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[1]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "bidir_dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 8;
defparam ram_block1a1.port_b_byte_enable_clock = "clock1";
defparam ram_block1a1.port_b_byte_enable_mask_width = 1;
defparam ram_block1a1.port_b_byte_size = 1;
defparam ram_block1a1.port_b_data_in_clock = "clock1";
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 255;
defparam ram_block1a1.port_b_logical_ram_depth = 256;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.port_b_write_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[2]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "bidir_dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 8;
defparam ram_block1a2.port_b_byte_enable_clock = "clock1";
defparam ram_block1a2.port_b_byte_enable_mask_width = 1;
defparam ram_block1a2.port_b_byte_size = 1;
defparam ram_block1a2.port_b_data_in_clock = "clock1";
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 255;
defparam ram_block1a2.port_b_logical_ram_depth = 256;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.port_b_write_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[3]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "bidir_dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 8;
defparam ram_block1a3.port_b_byte_enable_clock = "clock1";
defparam ram_block1a3.port_b_byte_enable_mask_width = 1;
defparam ram_block1a3.port_b_byte_size = 1;
defparam ram_block1a3.port_b_data_in_clock = "clock1";
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 255;
defparam ram_block1a3.port_b_logical_ram_depth = 256;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.port_b_write_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[4]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "bidir_dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 8;
defparam ram_block1a4.port_b_byte_enable_clock = "clock1";
defparam ram_block1a4.port_b_byte_enable_mask_width = 1;
defparam ram_block1a4.port_b_byte_size = 1;
defparam ram_block1a4.port_b_data_in_clock = "clock1";
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 255;
defparam ram_block1a4.port_b_logical_ram_depth = 256;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.port_b_write_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[5]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "bidir_dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 8;
defparam ram_block1a5.port_b_byte_enable_clock = "clock1";
defparam ram_block1a5.port_b_byte_enable_mask_width = 1;
defparam ram_block1a5.port_b_byte_size = 1;
defparam ram_block1a5.port_b_data_in_clock = "clock1";
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 255;
defparam ram_block1a5.port_b_logical_ram_depth = 256;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.port_b_write_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[6]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "bidir_dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 8;
defparam ram_block1a6.port_b_byte_enable_clock = "clock1";
defparam ram_block1a6.port_b_byte_enable_mask_width = 1;
defparam ram_block1a6.port_b_byte_size = 1;
defparam ram_block1a6.port_b_data_in_clock = "clock1";
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 255;
defparam ram_block1a6.port_b_logical_ram_depth = 256;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.port_b_write_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[7]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "bidir_dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 8;
defparam ram_block1a7.port_b_byte_enable_clock = "clock1";
defparam ram_block1a7.port_b_byte_enable_mask_width = 1;
defparam ram_block1a7.port_b_byte_size = 1;
defparam ram_block1a7.port_b_data_in_clock = "clock1";
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 255;
defparam ram_block1a7.port_b_logical_ram_depth = 256;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.port_b_write_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[8]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk1_core_clock_enable = "ena1";
defparam ram_block1a8.clk1_input_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "bidir_dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 8;
defparam ram_block1a8.port_b_byte_enable_clock = "clock1";
defparam ram_block1a8.port_b_byte_enable_mask_width = 1;
defparam ram_block1a8.port_b_byte_size = 1;
defparam ram_block1a8.port_b_data_in_clock = "clock1";
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 255;
defparam ram_block1a8.port_b_logical_ram_depth = 256;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.port_b_write_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[9]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk1_core_clock_enable = "ena1";
defparam ram_block1a9.clk1_input_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "bidir_dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 8;
defparam ram_block1a9.port_b_byte_enable_clock = "clock1";
defparam ram_block1a9.port_b_byte_enable_mask_width = 1;
defparam ram_block1a9.port_b_byte_size = 1;
defparam ram_block1a9.port_b_data_in_clock = "clock1";
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 255;
defparam ram_block1a9.port_b_logical_ram_depth = 256;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.port_b_write_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[10]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk1_core_clock_enable = "ena1";
defparam ram_block1a10.clk1_input_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "bidir_dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 8;
defparam ram_block1a10.port_b_byte_enable_clock = "clock1";
defparam ram_block1a10.port_b_byte_enable_mask_width = 1;
defparam ram_block1a10.port_b_byte_size = 1;
defparam ram_block1a10.port_b_data_in_clock = "clock1";
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 255;
defparam ram_block1a10.port_b_logical_ram_depth = 256;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.port_b_write_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[11]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk1_core_clock_enable = "ena1";
defparam ram_block1a11.clk1_input_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "bidir_dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 8;
defparam ram_block1a11.port_b_byte_enable_clock = "clock1";
defparam ram_block1a11.port_b_byte_enable_mask_width = 1;
defparam ram_block1a11.port_b_byte_size = 1;
defparam ram_block1a11.port_b_data_in_clock = "clock1";
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 255;
defparam ram_block1a11.port_b_logical_ram_depth = 256;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.port_b_write_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[12]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk1_core_clock_enable = "ena1";
defparam ram_block1a12.clk1_input_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "bidir_dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 8;
defparam ram_block1a12.port_b_byte_enable_clock = "clock1";
defparam ram_block1a12.port_b_byte_enable_mask_width = 1;
defparam ram_block1a12.port_b_byte_size = 1;
defparam ram_block1a12.port_b_data_in_clock = "clock1";
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 255;
defparam ram_block1a12.port_b_logical_ram_depth = 256;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.port_b_write_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[13]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk1_core_clock_enable = "ena1";
defparam ram_block1a13.clk1_input_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "bidir_dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 8;
defparam ram_block1a13.port_b_byte_enable_clock = "clock1";
defparam ram_block1a13.port_b_byte_enable_mask_width = 1;
defparam ram_block1a13.port_b_byte_size = 1;
defparam ram_block1a13.port_b_data_in_clock = "clock1";
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 255;
defparam ram_block1a13.port_b_logical_ram_depth = 256;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.port_b_write_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[14]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk1_core_clock_enable = "ena1";
defparam ram_block1a14.clk1_input_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "bidir_dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 8;
defparam ram_block1a14.port_b_byte_enable_clock = "clock1";
defparam ram_block1a14.port_b_byte_enable_mask_width = 1;
defparam ram_block1a14.port_b_byte_size = 1;
defparam ram_block1a14.port_b_data_in_clock = "clock1";
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 255;
defparam ram_block1a14.port_b_logical_ram_depth = 256;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.port_b_write_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[15]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk1_core_clock_enable = "ena1";
defparam ram_block1a15.clk1_input_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "bidir_dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 8;
defparam ram_block1a15.port_b_byte_enable_clock = "clock1";
defparam ram_block1a15.port_b_byte_enable_mask_width = 1;
defparam ram_block1a15.port_b_byte_size = 1;
defparam ram_block1a15.port_b_data_in_clock = "clock1";
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 255;
defparam ram_block1a15.port_b_logical_ram_depth = 256;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.port_b_write_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[16]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk1_core_clock_enable = "ena1";
defparam ram_block1a16.clk1_input_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "bidir_dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 8;
defparam ram_block1a16.port_b_byte_enable_clock = "clock1";
defparam ram_block1a16.port_b_byte_enable_mask_width = 1;
defparam ram_block1a16.port_b_byte_size = 1;
defparam ram_block1a16.port_b_data_in_clock = "clock1";
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 255;
defparam ram_block1a16.port_b_logical_ram_depth = 256;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.port_b_write_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[17]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk1_core_clock_enable = "ena1";
defparam ram_block1a17.clk1_input_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "bidir_dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 8;
defparam ram_block1a17.port_b_byte_enable_clock = "clock1";
defparam ram_block1a17.port_b_byte_enable_mask_width = 1;
defparam ram_block1a17.port_b_byte_size = 1;
defparam ram_block1a17.port_b_data_in_clock = "clock1";
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 255;
defparam ram_block1a17.port_b_logical_ram_depth = 256;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.port_b_write_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[18]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk1_core_clock_enable = "ena1";
defparam ram_block1a18.clk1_input_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "bidir_dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 8;
defparam ram_block1a18.port_b_byte_enable_clock = "clock1";
defparam ram_block1a18.port_b_byte_enable_mask_width = 1;
defparam ram_block1a18.port_b_byte_size = 1;
defparam ram_block1a18.port_b_data_in_clock = "clock1";
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 255;
defparam ram_block1a18.port_b_logical_ram_depth = 256;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.port_b_write_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[19]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk1_core_clock_enable = "ena1";
defparam ram_block1a19.clk1_input_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "bidir_dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 8;
defparam ram_block1a19.port_b_byte_enable_clock = "clock1";
defparam ram_block1a19.port_b_byte_enable_mask_width = 1;
defparam ram_block1a19.port_b_byte_size = 1;
defparam ram_block1a19.port_b_data_in_clock = "clock1";
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 255;
defparam ram_block1a19.port_b_logical_ram_depth = 256;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.port_b_write_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[20]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.clk1_core_clock_enable = "ena1";
defparam ram_block1a20.clk1_input_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "bidir_dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 8;
defparam ram_block1a20.port_b_byte_enable_clock = "clock1";
defparam ram_block1a20.port_b_byte_enable_mask_width = 1;
defparam ram_block1a20.port_b_byte_size = 1;
defparam ram_block1a20.port_b_data_in_clock = "clock1";
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 255;
defparam ram_block1a20.port_b_logical_ram_depth = 256;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.port_b_write_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[21]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.clk1_core_clock_enable = "ena1";
defparam ram_block1a21.clk1_input_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "bidir_dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 8;
defparam ram_block1a21.port_b_byte_enable_clock = "clock1";
defparam ram_block1a21.port_b_byte_enable_mask_width = 1;
defparam ram_block1a21.port_b_byte_size = 1;
defparam ram_block1a21.port_b_data_in_clock = "clock1";
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 255;
defparam ram_block1a21.port_b_logical_ram_depth = 256;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.port_b_write_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[22]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.clk1_core_clock_enable = "ena1";
defparam ram_block1a22.clk1_input_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "bidir_dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 8;
defparam ram_block1a22.port_b_byte_enable_clock = "clock1";
defparam ram_block1a22.port_b_byte_enable_mask_width = 1;
defparam ram_block1a22.port_b_byte_size = 1;
defparam ram_block1a22.port_b_data_in_clock = "clock1";
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 255;
defparam ram_block1a22.port_b_logical_ram_depth = 256;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.port_b_write_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[23]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.clk1_core_clock_enable = "ena1";
defparam ram_block1a23.clk1_input_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "bidir_dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 8;
defparam ram_block1a23.port_b_byte_enable_clock = "clock1";
defparam ram_block1a23.port_b_byte_enable_mask_width = 1;
defparam ram_block1a23.port_b_byte_size = 1;
defparam ram_block1a23.port_b_data_in_clock = "clock1";
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 255;
defparam ram_block1a23.port_b_logical_ram_depth = 256;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.port_b_write_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[24]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.clk1_core_clock_enable = "ena1";
defparam ram_block1a24.clk1_input_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "bidir_dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 8;
defparam ram_block1a24.port_b_byte_enable_clock = "clock1";
defparam ram_block1a24.port_b_byte_enable_mask_width = 1;
defparam ram_block1a24.port_b_byte_size = 1;
defparam ram_block1a24.port_b_data_in_clock = "clock1";
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 255;
defparam ram_block1a24.port_b_logical_ram_depth = 256;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.port_b_write_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[25]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.clk1_core_clock_enable = "ena1";
defparam ram_block1a25.clk1_input_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "bidir_dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 8;
defparam ram_block1a25.port_b_byte_enable_clock = "clock1";
defparam ram_block1a25.port_b_byte_enable_mask_width = 1;
defparam ram_block1a25.port_b_byte_size = 1;
defparam ram_block1a25.port_b_data_in_clock = "clock1";
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 255;
defparam ram_block1a25.port_b_logical_ram_depth = 256;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.port_b_write_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[26]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.clk1_core_clock_enable = "ena1";
defparam ram_block1a26.clk1_input_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "bidir_dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 8;
defparam ram_block1a26.port_b_byte_enable_clock = "clock1";
defparam ram_block1a26.port_b_byte_enable_mask_width = 1;
defparam ram_block1a26.port_b_byte_size = 1;
defparam ram_block1a26.port_b_data_in_clock = "clock1";
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 255;
defparam ram_block1a26.port_b_logical_ram_depth = 256;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.port_b_write_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[27]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.clk1_core_clock_enable = "ena1";
defparam ram_block1a27.clk1_input_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "bidir_dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 8;
defparam ram_block1a27.port_b_byte_enable_clock = "clock1";
defparam ram_block1a27.port_b_byte_enable_mask_width = 1;
defparam ram_block1a27.port_b_byte_size = 1;
defparam ram_block1a27.port_b_data_in_clock = "clock1";
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 255;
defparam ram_block1a27.port_b_logical_ram_depth = 256;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.port_b_write_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[28]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.clk1_core_clock_enable = "ena1";
defparam ram_block1a28.clk1_input_clock_enable = "ena1";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "bidir_dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 8;
defparam ram_block1a28.port_b_byte_enable_clock = "clock1";
defparam ram_block1a28.port_b_byte_enable_mask_width = 1;
defparam ram_block1a28.port_b_byte_size = 1;
defparam ram_block1a28.port_b_data_in_clock = "clock1";
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 255;
defparam ram_block1a28.port_b_logical_ram_depth = 256;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.port_b_write_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[29]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.clk1_core_clock_enable = "ena1";
defparam ram_block1a29.clk1_input_clock_enable = "ena1";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "bidir_dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 8;
defparam ram_block1a29.port_b_byte_enable_clock = "clock1";
defparam ram_block1a29.port_b_byte_enable_mask_width = 1;
defparam ram_block1a29.port_b_byte_size = 1;
defparam ram_block1a29.port_b_data_in_clock = "clock1";
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 255;
defparam ram_block1a29.port_b_logical_ram_depth = 256;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.port_b_write_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[30]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.clk1_core_clock_enable = "ena1";
defparam ram_block1a30.clk1_input_clock_enable = "ena1";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "bidir_dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 8;
defparam ram_block1a30.port_b_byte_enable_clock = "clock1";
defparam ram_block1a30.port_b_byte_enable_mask_width = 1;
defparam ram_block1a30.port_b_byte_size = 1;
defparam ram_block1a30.port_b_data_in_clock = "clock1";
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 255;
defparam ram_block1a30.port_b_logical_ram_depth = 256;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.port_b_write_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(!clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[31]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.clk1_core_clock_enable = "ena1";
defparam ram_block1a31.clk1_input_clock_enable = "ena1";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "Computer_System_Onchip_SRAM:onchip_sram|altsyncram:the_altsyncram|altsyncram_1k52:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "bidir_dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 8;
defparam ram_block1a31.port_b_byte_enable_clock = "clock1";
defparam ram_block1a31.port_b_byte_enable_mask_width = 1;
defparam ram_block1a31.port_b_byte_size = 1;
defparam ram_block1a31.port_b_data_in_clock = "clock1";
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 255;
defparam ram_block1a31.port_b_logical_ram_depth = 256;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.port_b_write_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

endmodule

module Computer_System_Computer_System_System_PLL (
	outclk_wire_1,
	outclk_wire_0,
	locked_wire_0,
	system_pll_ref_clk_clk,
	system_pll_ref_reset_reset)/* synthesis synthesis_greybox=0 */;
output 	outclk_wire_1;
output 	outclk_wire_0;
output 	locked_wire_0;
input 	system_pll_ref_clk_clk;
input 	system_pll_ref_reset_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_Computer_System_System_PLL_sys_pll sys_pll(
	.outclk_wire_1(outclk_wire_1),
	.outclk_wire_0(outclk_wire_0),
	.locked(locked_wire_0),
	.system_pll_ref_clk_clk(system_pll_ref_clk_clk),
	.system_pll_ref_reset_reset(system_pll_ref_reset_reset));

endmodule

module Computer_System_Computer_System_System_PLL_sys_pll (
	outclk_wire_1,
	outclk_wire_0,
	locked,
	system_pll_ref_clk_clk,
	system_pll_ref_reset_reset)/* synthesis synthesis_greybox=0 */;
output 	outclk_wire_1;
output 	outclk_wire_0;
output 	locked;
input 	system_pll_ref_clk_clk;
input 	system_pll_ref_reset_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



Computer_System_altera_pll_1 altera_pll_i(
	.outclk({outclk_wire_1,outclk_wire_0}),
	.locked(locked),
	.refclk(system_pll_ref_clk_clk),
	.rst(system_pll_ref_reset_reset));

endmodule

module Computer_System_altera_pll_1 (
	outclk,
	locked,
	refclk,
	rst)/* synthesis synthesis_greybox=0 */;
output 	[1:0] outclk;
output 	locked;
input 	refclk;
input 	rst;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fboutclk_wire[0] ;


generic_pll \general[1].gpll (
	.refclk(refclk),
	.fbclk(\fboutclk_wire[0] ),
	.rst(rst),
	.writerefclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writeoutclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writephaseshiftdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writedutycycledata(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.outclk(outclk[1]),
	.fboutclk(),
	.locked(),
	.readrefclkdata(),
	.readoutclkdata(),
	.readphaseshiftdata(),
	.readdutycycledata());
defparam \general[1].gpll .clock_name_global = "false";
defparam \general[1].gpll .duty_cycle = 50;
defparam \general[1].gpll .fractional_vco_multiplier = "false";
defparam \general[1].gpll .output_clock_frequency = "100.0 mhz";
defparam \general[1].gpll .phase_shift = "-3000 ps";
defparam \general[1].gpll .reference_clock_frequency = "50.0 mhz";
defparam \general[1].gpll .simulation_type = "timing";

generic_pll \general[0].gpll (
	.refclk(refclk),
	.fbclk(\fboutclk_wire[0] ),
	.rst(rst),
	.writerefclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writeoutclkdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writephaseshiftdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.writedutycycledata(64'b0000000000000000000000000000000000000000000000000000000000000000),
	.outclk(outclk[0]),
	.fboutclk(\fboutclk_wire[0] ),
	.locked(locked),
	.readrefclkdata(),
	.readoutclkdata(),
	.readphaseshiftdata(),
	.readdutycycledata());
defparam \general[0].gpll .clock_name_global = "false";
defparam \general[0].gpll .duty_cycle = 50;
defparam \general[0].gpll .fractional_vco_multiplier = "false";
defparam \general[0].gpll .output_clock_frequency = "100.0 mhz";
defparam \general[0].gpll .phase_shift = "0 ps";
defparam \general[0].gpll .reference_clock_frequency = "50.0 mhz";
defparam \general[0].gpll .simulation_type = "timing";

endmodule
